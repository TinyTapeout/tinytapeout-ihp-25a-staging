module tt_um_larva (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire clk_regs;
 wire bsq1r;
 wire \bsq[0] ;
 wire \bsq[10] ;
 wire \bsq[11] ;
 wire \bsq[12] ;
 wire \bsq[13] ;
 wire \bsq[14] ;
 wire \bsq[15] ;
 wire \bsq[16] ;
 wire \bsq[17] ;
 wire \bsq[18] ;
 wire \bsq[19] ;
 wire \bsq[1] ;
 wire \bsq[20] ;
 wire \bsq[21] ;
 wire \bsq[22] ;
 wire \bsq[23] ;
 wire \bsq[24] ;
 wire \bsq[25] ;
 wire \bsq[26] ;
 wire \bsq[27] ;
 wire \bsq[28] ;
 wire \bsq[29] ;
 wire \bsq[2] ;
 wire \bsq[3] ;
 wire \bsq[4] ;
 wire \bsq[5] ;
 wire \bsq[6] ;
 wire \bsq[7] ;
 wire \bsq[8] ;
 wire \bsq[9] ;
 wire cclk;
 wire \cdi[0] ;
 wire \cdi[10] ;
 wire \cdi[11] ;
 wire \cdi[12] ;
 wire \cdi[13] ;
 wire \cdi[14] ;
 wire \cdi[15] ;
 wire \cdi[16] ;
 wire \cdi[17] ;
 wire \cdi[18] ;
 wire \cdi[19] ;
 wire \cdi[1] ;
 wire \cdi[20] ;
 wire \cdi[21] ;
 wire \cdi[22] ;
 wire \cdi[23] ;
 wire \cdi[24] ;
 wire \cdi[25] ;
 wire \cdi[26] ;
 wire \cdi[27] ;
 wire \cdi[28] ;
 wire \cdi[29] ;
 wire \cdi[2] ;
 wire \cdi[30] ;
 wire \cdi[31] ;
 wire \cdi[3] ;
 wire \cdi[4] ;
 wire \cdi[5] ;
 wire \cdi[6] ;
 wire \cdi[7] ;
 wire \cdi[8] ;
 wire \cdi[9] ;
 wire \ckd[0] ;
 wire \ckd[1] ;
 wire \ckd[2] ;
 wire \cpu.Bimm[10] ;
 wire \cpu.Bimm[11] ;
 wire \cpu.Bimm[12] ;
 wire \cpu.Bimm[1] ;
 wire \cpu.Bimm[2] ;
 wire \cpu.Bimm[3] ;
 wire \cpu.Bimm[4] ;
 wire \cpu.Bimm[5] ;
 wire \cpu.Bimm[6] ;
 wire \cpu.Bimm[7] ;
 wire \cpu.Bimm[8] ;
 wire \cpu.Bimm[9] ;
 wire \cpu.IR[0] ;
 wire \cpu.IR[12] ;
 wire \cpu.IR[13] ;
 wire \cpu.IR[14] ;
 wire \cpu.IR[15] ;
 wire \cpu.IR[16] ;
 wire \cpu.IR[17] ;
 wire \cpu.IR[18] ;
 wire \cpu.IR[19] ;
 wire \cpu.IR[1] ;
 wire \cpu.IR[20] ;
 wire \cpu.IR[21] ;
 wire \cpu.IR[22] ;
 wire \cpu.IR[23] ;
 wire \cpu.IR[24] ;
 wire \cpu.IR[2] ;
 wire \cpu.IR[3] ;
 wire \cpu.IR[4] ;
 wire \cpu.IR[5] ;
 wire \cpu.IR[6] ;
 wire \cpu.PC[10] ;
 wire \cpu.PC[11] ;
 wire \cpu.PC[12] ;
 wire \cpu.PC[13] ;
 wire \cpu.PC[14] ;
 wire \cpu.PC[15] ;
 wire \cpu.PC[16] ;
 wire \cpu.PC[17] ;
 wire \cpu.PC[18] ;
 wire \cpu.PC[19] ;
 wire \cpu.PC[20] ;
 wire \cpu.PC[21] ;
 wire \cpu.PC[22] ;
 wire \cpu.PC[23] ;
 wire \cpu.PC[24] ;
 wire \cpu.PC[25] ;
 wire \cpu.PC[26] ;
 wire \cpu.PC[27] ;
 wire \cpu.PC[28] ;
 wire \cpu.PC[29] ;
 wire \cpu.PC[2] ;
 wire \cpu.PC[30] ;
 wire \cpu.PC[31] ;
 wire \cpu.PC[3] ;
 wire \cpu.PC[4] ;
 wire \cpu.PC[5] ;
 wire \cpu.PC[6] ;
 wire \cpu.PC[7] ;
 wire \cpu.PC[8] ;
 wire \cpu.PC[9] ;
 wire \cpu.PCci[10] ;
 wire \cpu.PCci[11] ;
 wire \cpu.PCci[12] ;
 wire \cpu.PCci[13] ;
 wire \cpu.PCci[14] ;
 wire \cpu.PCci[15] ;
 wire \cpu.PCci[16] ;
 wire \cpu.PCci[17] ;
 wire \cpu.PCci[18] ;
 wire \cpu.PCci[19] ;
 wire \cpu.PCci[20] ;
 wire \cpu.PCci[21] ;
 wire \cpu.PCci[22] ;
 wire \cpu.PCci[23] ;
 wire \cpu.PCci[24] ;
 wire \cpu.PCci[25] ;
 wire \cpu.PCci[26] ;
 wire \cpu.PCci[27] ;
 wire \cpu.PCci[28] ;
 wire \cpu.PCci[29] ;
 wire \cpu.PCci[2] ;
 wire \cpu.PCci[30] ;
 wire \cpu.PCci[31] ;
 wire \cpu.PCci[3] ;
 wire \cpu.PCci[4] ;
 wire \cpu.PCci[5] ;
 wire \cpu.PCci[6] ;
 wire \cpu.PCci[7] ;
 wire \cpu.PCci[8] ;
 wire \cpu.PCci[9] ;
 wire \cpu.PCreg0[10] ;
 wire \cpu.PCreg0[11] ;
 wire \cpu.PCreg0[12] ;
 wire \cpu.PCreg0[13] ;
 wire \cpu.PCreg0[14] ;
 wire \cpu.PCreg0[15] ;
 wire \cpu.PCreg0[16] ;
 wire \cpu.PCreg0[17] ;
 wire \cpu.PCreg0[18] ;
 wire \cpu.PCreg0[19] ;
 wire \cpu.PCreg0[20] ;
 wire \cpu.PCreg0[21] ;
 wire \cpu.PCreg0[22] ;
 wire \cpu.PCreg0[23] ;
 wire \cpu.PCreg0[24] ;
 wire \cpu.PCreg0[25] ;
 wire \cpu.PCreg0[26] ;
 wire \cpu.PCreg0[27] ;
 wire \cpu.PCreg0[28] ;
 wire \cpu.PCreg0[29] ;
 wire \cpu.PCreg0[2] ;
 wire \cpu.PCreg0[30] ;
 wire \cpu.PCreg0[31] ;
 wire \cpu.PCreg0[3] ;
 wire \cpu.PCreg0[4] ;
 wire \cpu.PCreg0[5] ;
 wire \cpu.PCreg0[6] ;
 wire \cpu.PCreg0[7] ;
 wire \cpu.PCreg0[8] ;
 wire \cpu.PCreg0[9] ;
 wire \cpu.PCreg1[10] ;
 wire \cpu.PCreg1[11] ;
 wire \cpu.PCreg1[12] ;
 wire \cpu.PCreg1[13] ;
 wire \cpu.PCreg1[14] ;
 wire \cpu.PCreg1[15] ;
 wire \cpu.PCreg1[16] ;
 wire \cpu.PCreg1[17] ;
 wire \cpu.PCreg1[18] ;
 wire \cpu.PCreg1[19] ;
 wire \cpu.PCreg1[20] ;
 wire \cpu.PCreg1[21] ;
 wire \cpu.PCreg1[22] ;
 wire \cpu.PCreg1[23] ;
 wire \cpu.PCreg1[24] ;
 wire \cpu.PCreg1[25] ;
 wire \cpu.PCreg1[26] ;
 wire \cpu.PCreg1[27] ;
 wire \cpu.PCreg1[28] ;
 wire \cpu.PCreg1[29] ;
 wire \cpu.PCreg1[2] ;
 wire \cpu.PCreg1[30] ;
 wire \cpu.PCreg1[31] ;
 wire \cpu.PCreg1[3] ;
 wire \cpu.PCreg1[4] ;
 wire \cpu.PCreg1[5] ;
 wire \cpu.PCreg1[6] ;
 wire \cpu.PCreg1[7] ;
 wire \cpu.PCreg1[8] ;
 wire \cpu.PCreg1[9] ;
 wire \cpu.mmode ;
 wire \cpu.opvalid ;
 wire \cpu.q0 ;
 wire \cpu.regs[10][0] ;
 wire \cpu.regs[10][10] ;
 wire \cpu.regs[10][11] ;
 wire \cpu.regs[10][12] ;
 wire \cpu.regs[10][13] ;
 wire \cpu.regs[10][14] ;
 wire \cpu.regs[10][15] ;
 wire \cpu.regs[10][16] ;
 wire \cpu.regs[10][17] ;
 wire \cpu.regs[10][18] ;
 wire \cpu.regs[10][19] ;
 wire \cpu.regs[10][1] ;
 wire \cpu.regs[10][20] ;
 wire \cpu.regs[10][21] ;
 wire \cpu.regs[10][22] ;
 wire \cpu.regs[10][23] ;
 wire \cpu.regs[10][24] ;
 wire \cpu.regs[10][25] ;
 wire \cpu.regs[10][26] ;
 wire \cpu.regs[10][27] ;
 wire \cpu.regs[10][28] ;
 wire \cpu.regs[10][29] ;
 wire \cpu.regs[10][2] ;
 wire \cpu.regs[10][30] ;
 wire \cpu.regs[10][31] ;
 wire \cpu.regs[10][3] ;
 wire \cpu.regs[10][4] ;
 wire \cpu.regs[10][5] ;
 wire \cpu.regs[10][6] ;
 wire \cpu.regs[10][7] ;
 wire \cpu.regs[10][8] ;
 wire \cpu.regs[10][9] ;
 wire \cpu.regs[11][0] ;
 wire \cpu.regs[11][10] ;
 wire \cpu.regs[11][11] ;
 wire \cpu.regs[11][12] ;
 wire \cpu.regs[11][13] ;
 wire \cpu.regs[11][14] ;
 wire \cpu.regs[11][15] ;
 wire \cpu.regs[11][16] ;
 wire \cpu.regs[11][17] ;
 wire \cpu.regs[11][18] ;
 wire \cpu.regs[11][19] ;
 wire \cpu.regs[11][1] ;
 wire \cpu.regs[11][20] ;
 wire \cpu.regs[11][21] ;
 wire \cpu.regs[11][22] ;
 wire \cpu.regs[11][23] ;
 wire \cpu.regs[11][24] ;
 wire \cpu.regs[11][25] ;
 wire \cpu.regs[11][26] ;
 wire \cpu.regs[11][27] ;
 wire \cpu.regs[11][28] ;
 wire \cpu.regs[11][29] ;
 wire \cpu.regs[11][2] ;
 wire \cpu.regs[11][30] ;
 wire \cpu.regs[11][31] ;
 wire \cpu.regs[11][3] ;
 wire \cpu.regs[11][4] ;
 wire \cpu.regs[11][5] ;
 wire \cpu.regs[11][6] ;
 wire \cpu.regs[11][7] ;
 wire \cpu.regs[11][8] ;
 wire \cpu.regs[11][9] ;
 wire \cpu.regs[12][0] ;
 wire \cpu.regs[12][10] ;
 wire \cpu.regs[12][11] ;
 wire \cpu.regs[12][12] ;
 wire \cpu.regs[12][13] ;
 wire \cpu.regs[12][14] ;
 wire \cpu.regs[12][15] ;
 wire \cpu.regs[12][16] ;
 wire \cpu.regs[12][17] ;
 wire \cpu.regs[12][18] ;
 wire \cpu.regs[12][19] ;
 wire \cpu.regs[12][1] ;
 wire \cpu.regs[12][20] ;
 wire \cpu.regs[12][21] ;
 wire \cpu.regs[12][22] ;
 wire \cpu.regs[12][23] ;
 wire \cpu.regs[12][24] ;
 wire \cpu.regs[12][25] ;
 wire \cpu.regs[12][26] ;
 wire \cpu.regs[12][27] ;
 wire \cpu.regs[12][28] ;
 wire \cpu.regs[12][29] ;
 wire \cpu.regs[12][2] ;
 wire \cpu.regs[12][30] ;
 wire \cpu.regs[12][31] ;
 wire \cpu.regs[12][3] ;
 wire \cpu.regs[12][4] ;
 wire \cpu.regs[12][5] ;
 wire \cpu.regs[12][6] ;
 wire \cpu.regs[12][7] ;
 wire \cpu.regs[12][8] ;
 wire \cpu.regs[12][9] ;
 wire \cpu.regs[13][0] ;
 wire \cpu.regs[13][10] ;
 wire \cpu.regs[13][11] ;
 wire \cpu.regs[13][12] ;
 wire \cpu.regs[13][13] ;
 wire \cpu.regs[13][14] ;
 wire \cpu.regs[13][15] ;
 wire \cpu.regs[13][16] ;
 wire \cpu.regs[13][17] ;
 wire \cpu.regs[13][18] ;
 wire \cpu.regs[13][19] ;
 wire \cpu.regs[13][1] ;
 wire \cpu.regs[13][20] ;
 wire \cpu.regs[13][21] ;
 wire \cpu.regs[13][22] ;
 wire \cpu.regs[13][23] ;
 wire \cpu.regs[13][24] ;
 wire \cpu.regs[13][25] ;
 wire \cpu.regs[13][26] ;
 wire \cpu.regs[13][27] ;
 wire \cpu.regs[13][28] ;
 wire \cpu.regs[13][29] ;
 wire \cpu.regs[13][2] ;
 wire \cpu.regs[13][30] ;
 wire \cpu.regs[13][31] ;
 wire \cpu.regs[13][3] ;
 wire \cpu.regs[13][4] ;
 wire \cpu.regs[13][5] ;
 wire \cpu.regs[13][6] ;
 wire \cpu.regs[13][7] ;
 wire \cpu.regs[13][8] ;
 wire \cpu.regs[13][9] ;
 wire \cpu.regs[14][0] ;
 wire \cpu.regs[14][10] ;
 wire \cpu.regs[14][11] ;
 wire \cpu.regs[14][12] ;
 wire \cpu.regs[14][13] ;
 wire \cpu.regs[14][14] ;
 wire \cpu.regs[14][15] ;
 wire \cpu.regs[14][16] ;
 wire \cpu.regs[14][17] ;
 wire \cpu.regs[14][18] ;
 wire \cpu.regs[14][19] ;
 wire \cpu.regs[14][1] ;
 wire \cpu.regs[14][20] ;
 wire \cpu.regs[14][21] ;
 wire \cpu.regs[14][22] ;
 wire \cpu.regs[14][23] ;
 wire \cpu.regs[14][24] ;
 wire \cpu.regs[14][25] ;
 wire \cpu.regs[14][26] ;
 wire \cpu.regs[14][27] ;
 wire \cpu.regs[14][28] ;
 wire \cpu.regs[14][29] ;
 wire \cpu.regs[14][2] ;
 wire \cpu.regs[14][30] ;
 wire \cpu.regs[14][31] ;
 wire \cpu.regs[14][3] ;
 wire \cpu.regs[14][4] ;
 wire \cpu.regs[14][5] ;
 wire \cpu.regs[14][6] ;
 wire \cpu.regs[14][7] ;
 wire \cpu.regs[14][8] ;
 wire \cpu.regs[14][9] ;
 wire \cpu.regs[15][0] ;
 wire \cpu.regs[15][10] ;
 wire \cpu.regs[15][11] ;
 wire \cpu.regs[15][12] ;
 wire \cpu.regs[15][13] ;
 wire \cpu.regs[15][14] ;
 wire \cpu.regs[15][15] ;
 wire \cpu.regs[15][16] ;
 wire \cpu.regs[15][17] ;
 wire \cpu.regs[15][18] ;
 wire \cpu.regs[15][19] ;
 wire \cpu.regs[15][1] ;
 wire \cpu.regs[15][20] ;
 wire \cpu.regs[15][21] ;
 wire \cpu.regs[15][22] ;
 wire \cpu.regs[15][23] ;
 wire \cpu.regs[15][24] ;
 wire \cpu.regs[15][25] ;
 wire \cpu.regs[15][26] ;
 wire \cpu.regs[15][27] ;
 wire \cpu.regs[15][28] ;
 wire \cpu.regs[15][29] ;
 wire \cpu.regs[15][2] ;
 wire \cpu.regs[15][30] ;
 wire \cpu.regs[15][31] ;
 wire \cpu.regs[15][3] ;
 wire \cpu.regs[15][4] ;
 wire \cpu.regs[15][5] ;
 wire \cpu.regs[15][6] ;
 wire \cpu.regs[15][7] ;
 wire \cpu.regs[15][8] ;
 wire \cpu.regs[15][9] ;
 wire \cpu.regs[1][0] ;
 wire \cpu.regs[1][10] ;
 wire \cpu.regs[1][11] ;
 wire \cpu.regs[1][12] ;
 wire \cpu.regs[1][13] ;
 wire \cpu.regs[1][14] ;
 wire \cpu.regs[1][15] ;
 wire \cpu.regs[1][16] ;
 wire \cpu.regs[1][17] ;
 wire \cpu.regs[1][18] ;
 wire \cpu.regs[1][19] ;
 wire \cpu.regs[1][1] ;
 wire \cpu.regs[1][20] ;
 wire \cpu.regs[1][21] ;
 wire \cpu.regs[1][22] ;
 wire \cpu.regs[1][23] ;
 wire \cpu.regs[1][24] ;
 wire \cpu.regs[1][25] ;
 wire \cpu.regs[1][26] ;
 wire \cpu.regs[1][27] ;
 wire \cpu.regs[1][28] ;
 wire \cpu.regs[1][29] ;
 wire \cpu.regs[1][2] ;
 wire \cpu.regs[1][30] ;
 wire \cpu.regs[1][31] ;
 wire \cpu.regs[1][3] ;
 wire \cpu.regs[1][4] ;
 wire \cpu.regs[1][5] ;
 wire \cpu.regs[1][6] ;
 wire \cpu.regs[1][7] ;
 wire \cpu.regs[1][8] ;
 wire \cpu.regs[1][9] ;
 wire \cpu.regs[2][0] ;
 wire \cpu.regs[2][10] ;
 wire \cpu.regs[2][11] ;
 wire \cpu.regs[2][12] ;
 wire \cpu.regs[2][13] ;
 wire \cpu.regs[2][14] ;
 wire \cpu.regs[2][15] ;
 wire \cpu.regs[2][16] ;
 wire \cpu.regs[2][17] ;
 wire \cpu.regs[2][18] ;
 wire \cpu.regs[2][19] ;
 wire \cpu.regs[2][1] ;
 wire \cpu.regs[2][20] ;
 wire \cpu.regs[2][21] ;
 wire \cpu.regs[2][22] ;
 wire \cpu.regs[2][23] ;
 wire \cpu.regs[2][24] ;
 wire \cpu.regs[2][25] ;
 wire \cpu.regs[2][26] ;
 wire \cpu.regs[2][27] ;
 wire \cpu.regs[2][28] ;
 wire \cpu.regs[2][29] ;
 wire \cpu.regs[2][2] ;
 wire \cpu.regs[2][30] ;
 wire \cpu.regs[2][31] ;
 wire \cpu.regs[2][3] ;
 wire \cpu.regs[2][4] ;
 wire \cpu.regs[2][5] ;
 wire \cpu.regs[2][6] ;
 wire \cpu.regs[2][7] ;
 wire \cpu.regs[2][8] ;
 wire \cpu.regs[2][9] ;
 wire \cpu.regs[3][0] ;
 wire \cpu.regs[3][10] ;
 wire \cpu.regs[3][11] ;
 wire \cpu.regs[3][12] ;
 wire \cpu.regs[3][13] ;
 wire \cpu.regs[3][14] ;
 wire \cpu.regs[3][15] ;
 wire \cpu.regs[3][16] ;
 wire \cpu.regs[3][17] ;
 wire \cpu.regs[3][18] ;
 wire \cpu.regs[3][19] ;
 wire \cpu.regs[3][1] ;
 wire \cpu.regs[3][20] ;
 wire \cpu.regs[3][21] ;
 wire \cpu.regs[3][22] ;
 wire \cpu.regs[3][23] ;
 wire \cpu.regs[3][24] ;
 wire \cpu.regs[3][25] ;
 wire \cpu.regs[3][26] ;
 wire \cpu.regs[3][27] ;
 wire \cpu.regs[3][28] ;
 wire \cpu.regs[3][29] ;
 wire \cpu.regs[3][2] ;
 wire \cpu.regs[3][30] ;
 wire \cpu.regs[3][31] ;
 wire \cpu.regs[3][3] ;
 wire \cpu.regs[3][4] ;
 wire \cpu.regs[3][5] ;
 wire \cpu.regs[3][6] ;
 wire \cpu.regs[3][7] ;
 wire \cpu.regs[3][8] ;
 wire \cpu.regs[3][9] ;
 wire \cpu.regs[4][0] ;
 wire \cpu.regs[4][10] ;
 wire \cpu.regs[4][11] ;
 wire \cpu.regs[4][12] ;
 wire \cpu.regs[4][13] ;
 wire \cpu.regs[4][14] ;
 wire \cpu.regs[4][15] ;
 wire \cpu.regs[4][16] ;
 wire \cpu.regs[4][17] ;
 wire \cpu.regs[4][18] ;
 wire \cpu.regs[4][19] ;
 wire \cpu.regs[4][1] ;
 wire \cpu.regs[4][20] ;
 wire \cpu.regs[4][21] ;
 wire \cpu.regs[4][22] ;
 wire \cpu.regs[4][23] ;
 wire \cpu.regs[4][24] ;
 wire \cpu.regs[4][25] ;
 wire \cpu.regs[4][26] ;
 wire \cpu.regs[4][27] ;
 wire \cpu.regs[4][28] ;
 wire \cpu.regs[4][29] ;
 wire \cpu.regs[4][2] ;
 wire \cpu.regs[4][30] ;
 wire \cpu.regs[4][31] ;
 wire \cpu.regs[4][3] ;
 wire \cpu.regs[4][4] ;
 wire \cpu.regs[4][5] ;
 wire \cpu.regs[4][6] ;
 wire \cpu.regs[4][7] ;
 wire \cpu.regs[4][8] ;
 wire \cpu.regs[4][9] ;
 wire \cpu.regs[5][0] ;
 wire \cpu.regs[5][10] ;
 wire \cpu.regs[5][11] ;
 wire \cpu.regs[5][12] ;
 wire \cpu.regs[5][13] ;
 wire \cpu.regs[5][14] ;
 wire \cpu.regs[5][15] ;
 wire \cpu.regs[5][16] ;
 wire \cpu.regs[5][17] ;
 wire \cpu.regs[5][18] ;
 wire \cpu.regs[5][19] ;
 wire \cpu.regs[5][1] ;
 wire \cpu.regs[5][20] ;
 wire \cpu.regs[5][21] ;
 wire \cpu.regs[5][22] ;
 wire \cpu.regs[5][23] ;
 wire \cpu.regs[5][24] ;
 wire \cpu.regs[5][25] ;
 wire \cpu.regs[5][26] ;
 wire \cpu.regs[5][27] ;
 wire \cpu.regs[5][28] ;
 wire \cpu.regs[5][29] ;
 wire \cpu.regs[5][2] ;
 wire \cpu.regs[5][30] ;
 wire \cpu.regs[5][31] ;
 wire \cpu.regs[5][3] ;
 wire \cpu.regs[5][4] ;
 wire \cpu.regs[5][5] ;
 wire \cpu.regs[5][6] ;
 wire \cpu.regs[5][7] ;
 wire \cpu.regs[5][8] ;
 wire \cpu.regs[5][9] ;
 wire \cpu.regs[6][0] ;
 wire \cpu.regs[6][10] ;
 wire \cpu.regs[6][11] ;
 wire \cpu.regs[6][12] ;
 wire \cpu.regs[6][13] ;
 wire \cpu.regs[6][14] ;
 wire \cpu.regs[6][15] ;
 wire \cpu.regs[6][16] ;
 wire \cpu.regs[6][17] ;
 wire \cpu.regs[6][18] ;
 wire \cpu.regs[6][19] ;
 wire \cpu.regs[6][1] ;
 wire \cpu.regs[6][20] ;
 wire \cpu.regs[6][21] ;
 wire \cpu.regs[6][22] ;
 wire \cpu.regs[6][23] ;
 wire \cpu.regs[6][24] ;
 wire \cpu.regs[6][25] ;
 wire \cpu.regs[6][26] ;
 wire \cpu.regs[6][27] ;
 wire \cpu.regs[6][28] ;
 wire \cpu.regs[6][29] ;
 wire \cpu.regs[6][2] ;
 wire \cpu.regs[6][30] ;
 wire \cpu.regs[6][31] ;
 wire \cpu.regs[6][3] ;
 wire \cpu.regs[6][4] ;
 wire \cpu.regs[6][5] ;
 wire \cpu.regs[6][6] ;
 wire \cpu.regs[6][7] ;
 wire \cpu.regs[6][8] ;
 wire \cpu.regs[6][9] ;
 wire \cpu.regs[7][0] ;
 wire \cpu.regs[7][10] ;
 wire \cpu.regs[7][11] ;
 wire \cpu.regs[7][12] ;
 wire \cpu.regs[7][13] ;
 wire \cpu.regs[7][14] ;
 wire \cpu.regs[7][15] ;
 wire \cpu.regs[7][16] ;
 wire \cpu.regs[7][17] ;
 wire \cpu.regs[7][18] ;
 wire \cpu.regs[7][19] ;
 wire \cpu.regs[7][1] ;
 wire \cpu.regs[7][20] ;
 wire \cpu.regs[7][21] ;
 wire \cpu.regs[7][22] ;
 wire \cpu.regs[7][23] ;
 wire \cpu.regs[7][24] ;
 wire \cpu.regs[7][25] ;
 wire \cpu.regs[7][26] ;
 wire \cpu.regs[7][27] ;
 wire \cpu.regs[7][28] ;
 wire \cpu.regs[7][29] ;
 wire \cpu.regs[7][2] ;
 wire \cpu.regs[7][30] ;
 wire \cpu.regs[7][31] ;
 wire \cpu.regs[7][3] ;
 wire \cpu.regs[7][4] ;
 wire \cpu.regs[7][5] ;
 wire \cpu.regs[7][6] ;
 wire \cpu.regs[7][7] ;
 wire \cpu.regs[7][8] ;
 wire \cpu.regs[7][9] ;
 wire \cpu.regs[8][0] ;
 wire \cpu.regs[8][10] ;
 wire \cpu.regs[8][11] ;
 wire \cpu.regs[8][12] ;
 wire \cpu.regs[8][13] ;
 wire \cpu.regs[8][14] ;
 wire \cpu.regs[8][15] ;
 wire \cpu.regs[8][16] ;
 wire \cpu.regs[8][17] ;
 wire \cpu.regs[8][18] ;
 wire \cpu.regs[8][19] ;
 wire \cpu.regs[8][1] ;
 wire \cpu.regs[8][20] ;
 wire \cpu.regs[8][21] ;
 wire \cpu.regs[8][22] ;
 wire \cpu.regs[8][23] ;
 wire \cpu.regs[8][24] ;
 wire \cpu.regs[8][25] ;
 wire \cpu.regs[8][26] ;
 wire \cpu.regs[8][27] ;
 wire \cpu.regs[8][28] ;
 wire \cpu.regs[8][29] ;
 wire \cpu.regs[8][2] ;
 wire \cpu.regs[8][30] ;
 wire \cpu.regs[8][31] ;
 wire \cpu.regs[8][3] ;
 wire \cpu.regs[8][4] ;
 wire \cpu.regs[8][5] ;
 wire \cpu.regs[8][6] ;
 wire \cpu.regs[8][7] ;
 wire \cpu.regs[8][8] ;
 wire \cpu.regs[8][9] ;
 wire \cpu.regs[9][0] ;
 wire \cpu.regs[9][10] ;
 wire \cpu.regs[9][11] ;
 wire \cpu.regs[9][12] ;
 wire \cpu.regs[9][13] ;
 wire \cpu.regs[9][14] ;
 wire \cpu.regs[9][15] ;
 wire \cpu.regs[9][16] ;
 wire \cpu.regs[9][17] ;
 wire \cpu.regs[9][18] ;
 wire \cpu.regs[9][19] ;
 wire \cpu.regs[9][1] ;
 wire \cpu.regs[9][20] ;
 wire \cpu.regs[9][21] ;
 wire \cpu.regs[9][22] ;
 wire \cpu.regs[9][23] ;
 wire \cpu.regs[9][24] ;
 wire \cpu.regs[9][25] ;
 wire \cpu.regs[9][26] ;
 wire \cpu.regs[9][27] ;
 wire \cpu.regs[9][28] ;
 wire \cpu.regs[9][29] ;
 wire \cpu.regs[9][2] ;
 wire \cpu.regs[9][30] ;
 wire \cpu.regs[9][31] ;
 wire \cpu.regs[9][3] ;
 wire \cpu.regs[9][4] ;
 wire \cpu.regs[9][5] ;
 wire \cpu.regs[9][6] ;
 wire \cpu.regs[9][7] ;
 wire \cpu.regs[9][8] ;
 wire \cpu.regs[9][9] ;
 wire exintest;
 wire \irqen[0] ;
 wire \irqen[1] ;
 wire \irqen[2] ;
 wire \irqen[3] ;
 wire \irqen[4] ;
 wire \irqvect[0][0] ;
 wire \irqvect[0][10] ;
 wire \irqvect[0][11] ;
 wire \irqvect[0][12] ;
 wire \irqvect[0][13] ;
 wire \irqvect[0][14] ;
 wire \irqvect[0][15] ;
 wire \irqvect[0][16] ;
 wire \irqvect[0][17] ;
 wire \irqvect[0][18] ;
 wire \irqvect[0][19] ;
 wire \irqvect[0][1] ;
 wire \irqvect[0][20] ;
 wire \irqvect[0][21] ;
 wire \irqvect[0][22] ;
 wire \irqvect[0][23] ;
 wire \irqvect[0][24] ;
 wire \irqvect[0][25] ;
 wire \irqvect[0][26] ;
 wire \irqvect[0][27] ;
 wire \irqvect[0][28] ;
 wire \irqvect[0][29] ;
 wire \irqvect[0][2] ;
 wire \irqvect[0][3] ;
 wire \irqvect[0][4] ;
 wire \irqvect[0][5] ;
 wire \irqvect[0][6] ;
 wire \irqvect[0][7] ;
 wire \irqvect[0][8] ;
 wire \irqvect[0][9] ;
 wire \irqvect[1][0] ;
 wire \irqvect[1][10] ;
 wire \irqvect[1][11] ;
 wire \irqvect[1][12] ;
 wire \irqvect[1][13] ;
 wire \irqvect[1][14] ;
 wire \irqvect[1][15] ;
 wire \irqvect[1][16] ;
 wire \irqvect[1][17] ;
 wire \irqvect[1][18] ;
 wire \irqvect[1][19] ;
 wire \irqvect[1][1] ;
 wire \irqvect[1][20] ;
 wire \irqvect[1][21] ;
 wire \irqvect[1][22] ;
 wire \irqvect[1][23] ;
 wire \irqvect[1][24] ;
 wire \irqvect[1][25] ;
 wire \irqvect[1][26] ;
 wire \irqvect[1][27] ;
 wire \irqvect[1][28] ;
 wire \irqvect[1][29] ;
 wire \irqvect[1][2] ;
 wire \irqvect[1][3] ;
 wire \irqvect[1][4] ;
 wire \irqvect[1][5] ;
 wire \irqvect[1][6] ;
 wire \irqvect[1][7] ;
 wire \irqvect[1][8] ;
 wire \irqvect[1][9] ;
 wire \irqvect[2][0] ;
 wire \irqvect[2][10] ;
 wire \irqvect[2][11] ;
 wire \irqvect[2][12] ;
 wire \irqvect[2][13] ;
 wire \irqvect[2][14] ;
 wire \irqvect[2][15] ;
 wire \irqvect[2][16] ;
 wire \irqvect[2][17] ;
 wire \irqvect[2][18] ;
 wire \irqvect[2][19] ;
 wire \irqvect[2][1] ;
 wire \irqvect[2][20] ;
 wire \irqvect[2][21] ;
 wire \irqvect[2][22] ;
 wire \irqvect[2][23] ;
 wire \irqvect[2][24] ;
 wire \irqvect[2][25] ;
 wire \irqvect[2][26] ;
 wire \irqvect[2][27] ;
 wire \irqvect[2][28] ;
 wire \irqvect[2][29] ;
 wire \irqvect[2][2] ;
 wire \irqvect[2][3] ;
 wire \irqvect[2][4] ;
 wire \irqvect[2][5] ;
 wire \irqvect[2][6] ;
 wire \irqvect[2][7] ;
 wire \irqvect[2][8] ;
 wire \irqvect[2][9] ;
 wire \irqvect[3][0] ;
 wire \irqvect[3][10] ;
 wire \irqvect[3][11] ;
 wire \irqvect[3][12] ;
 wire \irqvect[3][13] ;
 wire \irqvect[3][14] ;
 wire \irqvect[3][15] ;
 wire \irqvect[3][16] ;
 wire \irqvect[3][17] ;
 wire \irqvect[3][18] ;
 wire \irqvect[3][19] ;
 wire \irqvect[3][1] ;
 wire \irqvect[3][20] ;
 wire \irqvect[3][21] ;
 wire \irqvect[3][22] ;
 wire \irqvect[3][23] ;
 wire \irqvect[3][24] ;
 wire \irqvect[3][25] ;
 wire \irqvect[3][26] ;
 wire \irqvect[3][27] ;
 wire \irqvect[3][28] ;
 wire \irqvect[3][29] ;
 wire \irqvect[3][2] ;
 wire \irqvect[3][3] ;
 wire \irqvect[3][4] ;
 wire \irqvect[3][5] ;
 wire \irqvect[3][6] ;
 wire \irqvect[3][7] ;
 wire \irqvect[3][8] ;
 wire \irqvect[3][9] ;
 wire jclk;
 wire \jtag0.bssh[0] ;
 wire \jtag0.bssh[10] ;
 wire \jtag0.bssh[11] ;
 wire \jtag0.bssh[12] ;
 wire \jtag0.bssh[13] ;
 wire \jtag0.bssh[14] ;
 wire \jtag0.bssh[15] ;
 wire \jtag0.bssh[16] ;
 wire \jtag0.bssh[17] ;
 wire \jtag0.bssh[18] ;
 wire \jtag0.bssh[19] ;
 wire \jtag0.bssh[1] ;
 wire \jtag0.bssh[20] ;
 wire \jtag0.bssh[21] ;
 wire \jtag0.bssh[22] ;
 wire \jtag0.bssh[23] ;
 wire \jtag0.bssh[24] ;
 wire \jtag0.bssh[25] ;
 wire \jtag0.bssh[26] ;
 wire \jtag0.bssh[27] ;
 wire \jtag0.bssh[28] ;
 wire \jtag0.bssh[29] ;
 wire \jtag0.bssh[2] ;
 wire \jtag0.bssh[3] ;
 wire \jtag0.bssh[4] ;
 wire \jtag0.bssh[5] ;
 wire \jtag0.bssh[6] ;
 wire \jtag0.bssh[7] ;
 wire \jtag0.bssh[8] ;
 wire \jtag0.bssh[9] ;
 wire \jtag0.byp ;
 wire \jtag0.idr[0] ;
 wire \jtag0.idr[10] ;
 wire \jtag0.idr[11] ;
 wire \jtag0.idr[12] ;
 wire \jtag0.idr[13] ;
 wire \jtag0.idr[14] ;
 wire \jtag0.idr[15] ;
 wire \jtag0.idr[16] ;
 wire \jtag0.idr[17] ;
 wire \jtag0.idr[18] ;
 wire \jtag0.idr[19] ;
 wire \jtag0.idr[1] ;
 wire \jtag0.idr[20] ;
 wire \jtag0.idr[21] ;
 wire \jtag0.idr[22] ;
 wire \jtag0.idr[23] ;
 wire \jtag0.idr[24] ;
 wire \jtag0.idr[25] ;
 wire \jtag0.idr[26] ;
 wire \jtag0.idr[27] ;
 wire \jtag0.idr[28] ;
 wire \jtag0.idr[29] ;
 wire \jtag0.idr[2] ;
 wire \jtag0.idr[30] ;
 wire \jtag0.idr[31] ;
 wire \jtag0.idr[3] ;
 wire \jtag0.idr[4] ;
 wire \jtag0.idr[5] ;
 wire \jtag0.idr[6] ;
 wire \jtag0.idr[7] ;
 wire \jtag0.idr[8] ;
 wire \jtag0.idr[9] ;
 wire \jtag0.ir[0] ;
 wire \jtag0.ir[1] ;
 wire \jtag0.ir[2] ;
 wire \jtag0.irsh[0] ;
 wire \jtag0.irsh[1] ;
 wire \jtag0.irsh[2] ;
 wire \jtag0.stdi ;
 wire \jtag0.stms ;
 wire \jtag0.tapst[0] ;
 wire \jtag0.tapst[1] ;
 wire \jtag0.tapst[2] ;
 wire \jtag0.tapst[3] ;
 wire \pwm[0] ;
 wire \pwm[1] ;
 wire \pwm[2] ;
 wire \pwm[3] ;
 wire \pwm[4] ;
 wire \pwm[5] ;
 wire \pwm[6] ;
 wire \pwm[7] ;
 wire \pwmbuf[0] ;
 wire \pwmbuf[1] ;
 wire \pwmbuf[2] ;
 wire \pwmbuf[3] ;
 wire \pwmbuf[4] ;
 wire \pwmbuf[5] ;
 wire \pwmbuf[6] ;
 wire \pwmbuf[7] ;
 wire \pwmc[0] ;
 wire \pwmc[1] ;
 wire \pwmc[2] ;
 wire \pwmc[3] ;
 wire \pwmc[4] ;
 wire \pwmc[5] ;
 wire \pwmc[6] ;
 wire \pwmc[7] ;
 wire pwmirq;
 wire pwmout;
 wire pwmpin;
 wire rxd;
 wire \tcount[0] ;
 wire \tcount[10] ;
 wire \tcount[11] ;
 wire \tcount[12] ;
 wire \tcount[13] ;
 wire \tcount[14] ;
 wire \tcount[15] ;
 wire \tcount[16] ;
 wire \tcount[17] ;
 wire \tcount[18] ;
 wire \tcount[19] ;
 wire \tcount[1] ;
 wire \tcount[20] ;
 wire \tcount[21] ;
 wire \tcount[22] ;
 wire \tcount[23] ;
 wire \tcount[24] ;
 wire \tcount[25] ;
 wire \tcount[26] ;
 wire \tcount[27] ;
 wire \tcount[28] ;
 wire \tcount[29] ;
 wire \tcount[2] ;
 wire \tcount[30] ;
 wire \tcount[31] ;
 wire \tcount[3] ;
 wire \tcount[4] ;
 wire \tcount[5] ;
 wire \tcount[6] ;
 wire \tcount[7] ;
 wire \tcount[8] ;
 wire \tcount[9] ;
 wire txd;
 wire \uart0.q[0] ;
 wire \uart0.q[1] ;
 wire \uart0.q[2] ;
 wire \uart0.q[3] ;
 wire \uart0.q[4] ;
 wire \uart0.q[5] ;
 wire \uart0.q[6] ;
 wire \uart0.q[7] ;
 wire \uart0.rxdiv[0] ;
 wire \uart0.rxdiv[1] ;
 wire \uart0.rxdiv[2] ;
 wire \uart0.rxdiv[3] ;
 wire \uart0.rxdiv[4] ;
 wire \uart0.rxdiv[5] ;
 wire \uart0.rxoverr ;
 wire \uart0.rxreg[0] ;
 wire \uart0.rxreg[1] ;
 wire \uart0.rxvalid ;
 wire \uart0.txbitcnt[0] ;
 wire \uart0.txbitcnt[1] ;
 wire \uart0.txbitcnt[2] ;
 wire \uart0.txbitcnt[3] ;
 wire \uart0.txdiv[0] ;
 wire \uart0.txdiv[1] ;
 wire \uart0.txdiv[2] ;
 wire \uart0.txdiv[3] ;
 wire \uart0.txdiv[4] ;
 wire \uart0.txdiv[5] ;
 wire \uart0.txsh[1] ;
 wire \uart0.txsh[2] ;
 wire \uart0.txsh[3] ;
 wire \uart0.txsh[4] ;
 wire \uart0.txsh[5] ;
 wire \uart0.txsh[6] ;
 wire \uart0.txsh[7] ;
 wire \uart0.txsh[8] ;
 wire \uart0.urxbuffer[8] ;
 wire \uart0.urxsh[0] ;
 wire \uart0.urxsh[1] ;
 wire \uart0.urxsh[2] ;
 wire \uart0.urxsh[3] ;
 wire \uart0.urxsh[4] ;
 wire \uart0.urxsh[5] ;
 wire \uart0.urxsh[6] ;
 wire \uart0.urxsh[7] ;
 wire \uart0.urxsh[8] ;
 wire \uart0.urxsh[9] ;
 wire udirty;
 wire \xdi[0] ;
 wire \xdi[10] ;
 wire \xdi[11] ;
 wire \xdi[12] ;
 wire \xdi[13] ;
 wire \xdi[14] ;
 wire \xdi[15] ;
 wire \xdi[16] ;
 wire \xdi[17] ;
 wire \xdi[18] ;
 wire \xdi[19] ;
 wire \xdi[1] ;
 wire \xdi[20] ;
 wire \xdi[21] ;
 wire \xdi[22] ;
 wire \xdi[23] ;
 wire \xdi[2] ;
 wire \xdi[3] ;
 wire \xdi[4] ;
 wire \xdi[5] ;
 wire \xdi[6] ;
 wire \xdi[7] ;
 wire \xdi[8] ;
 wire \xdi[9] ;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire jclk_regs;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire clknet_0_jclk;
 wire clknet_1_0__leaf_jclk;
 wire clknet_1_1__leaf_jclk;
 wire clknet_0_jclk_regs;
 wire clknet_2_0__leaf_jclk_regs;
 wire clknet_2_1__leaf_jclk_regs;
 wire clknet_2_2__leaf_jclk_regs;
 wire clknet_2_3__leaf_jclk_regs;
 wire clknet_0__02583_;
 wire clknet_1_0__leaf__02583_;
 wire clknet_1_1__leaf__02583_;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire delaynet_2_clk;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;

 sg13g2_inv_1 _06951_ (.Y(_01539_),
    .A(\jtag0.irsh[0] ));
 sg13g2_inv_1 _06952_ (.Y(_01540_),
    .A(\uart0.rxvalid ));
 sg13g2_inv_1 _06953_ (.Y(_01541_),
    .A(\uart0.q[2] ));
 sg13g2_inv_1 _06954_ (.Y(_01542_),
    .A(\uart0.txbitcnt[2] ));
 sg13g2_inv_1 _06955_ (.Y(_01543_),
    .A(\jtag0.bssh[29] ));
 sg13g2_inv_1 _06956_ (.Y(_01544_),
    .A(\jtag0.bssh[28] ));
 sg13g2_inv_1 _06957_ (.Y(_01545_),
    .A(\jtag0.bssh[27] ));
 sg13g2_inv_1 _06958_ (.Y(_01546_),
    .A(\jtag0.bssh[24] ));
 sg13g2_inv_1 _06959_ (.Y(_01547_),
    .A(\jtag0.bssh[23] ));
 sg13g2_inv_1 _06960_ (.Y(_01548_),
    .A(\jtag0.bssh[22] ));
 sg13g2_inv_1 _06961_ (.Y(_01549_),
    .A(\jtag0.bssh[21] ));
 sg13g2_inv_1 _06962_ (.Y(_01550_),
    .A(\jtag0.bssh[18] ));
 sg13g2_inv_1 _06963_ (.Y(_01551_),
    .A(\jtag0.bssh[17] ));
 sg13g2_inv_1 _06964_ (.Y(_01552_),
    .A(\jtag0.bssh[16] ));
 sg13g2_inv_1 _06965_ (.Y(_01553_),
    .A(\jtag0.bssh[15] ));
 sg13g2_inv_1 _06966_ (.Y(_01554_),
    .A(\jtag0.bssh[0] ));
 sg13g2_inv_1 _06967_ (.Y(_01555_),
    .A(\jtag0.idr[19] ));
 sg13g2_inv_1 _06968_ (.Y(_01556_),
    .A(\jtag0.idr[18] ));
 sg13g2_inv_1 _06969_ (.Y(_01557_),
    .A(\jtag0.idr[15] ));
 sg13g2_inv_1 _06970_ (.Y(_01558_),
    .A(\jtag0.idr[14] ));
 sg13g2_inv_1 _06971_ (.Y(_01559_),
    .A(\jtag0.idr[13] ));
 sg13g2_inv_1 _06972_ (.Y(_01560_),
    .A(\jtag0.idr[12] ));
 sg13g2_inv_1 _06973_ (.Y(_01561_),
    .A(\jtag0.idr[11] ));
 sg13g2_inv_1 _06974_ (.Y(_01562_),
    .A(\jtag0.idr[10] ));
 sg13g2_inv_1 _06975_ (.Y(_01563_),
    .A(\jtag0.idr[9] ));
 sg13g2_inv_1 _06976_ (.Y(_01564_),
    .A(\jtag0.idr[8] ));
 sg13g2_inv_1 _06977_ (.Y(_01565_),
    .A(\jtag0.idr[7] ));
 sg13g2_inv_1 _06978_ (.Y(_01566_),
    .A(\jtag0.idr[6] ));
 sg13g2_inv_1 _06979_ (.Y(_01567_),
    .A(\jtag0.idr[5] ));
 sg13g2_inv_1 _06980_ (.Y(_01568_),
    .A(\jtag0.idr[4] ));
 sg13g2_inv_1 _06981_ (.Y(_01569_),
    .A(\jtag0.idr[3] ));
 sg13g2_inv_1 _06982_ (.Y(_01570_),
    .A(\jtag0.idr[2] ));
 sg13g2_inv_1 _06983_ (.Y(_01571_),
    .A(\jtag0.idr[1] ));
 sg13g2_inv_1 _06984_ (.Y(_01572_),
    .A(\jtag0.idr[0] ));
 sg13g2_inv_1 _06985_ (.Y(_01573_),
    .A(\jtag0.ir[0] ));
 sg13g2_inv_1 _06986_ (.Y(_01574_),
    .A(_00572_));
 sg13g2_inv_1 _06987_ (.Y(_01575_),
    .A(net3638));
 sg13g2_inv_1 _06988_ (.Y(_01576_),
    .A(_00200_));
 sg13g2_inv_1 _06989_ (.Y(_01577_),
    .A(_00456_));
 sg13g2_inv_1 _06990_ (.Y(_01578_),
    .A(_00328_));
 sg13g2_inv_1 _06991_ (.Y(_01579_),
    .A(_00520_));
 sg13g2_inv_1 _06992_ (.Y(_01580_),
    .A(_00201_));
 sg13g2_inv_1 _06993_ (.Y(_01581_),
    .A(_00425_));
 sg13g2_inv_1 _06994_ (.Y(_01582_),
    .A(_00202_));
 sg13g2_inv_1 _06995_ (.Y(_01583_),
    .A(_00458_));
 sg13g2_inv_1 _06996_ (.Y(_01584_),
    .A(_00330_));
 sg13g2_inv_1 _06997_ (.Y(_01585_),
    .A(_00522_));
 sg13g2_inv_1 _06998_ (.Y(_01586_),
    .A(_00426_));
 sg13g2_inv_1 _06999_ (.Y(_01587_),
    .A(_00203_));
 sg13g2_inv_1 _07000_ (.Y(_01588_),
    .A(_00459_));
 sg13g2_inv_1 _07001_ (.Y(_01589_),
    .A(_00331_));
 sg13g2_inv_1 _07002_ (.Y(_01590_),
    .A(_00427_));
 sg13g2_inv_1 _07003_ (.Y(_01591_),
    .A(_00204_));
 sg13g2_inv_1 _07004_ (.Y(_01592_),
    .A(_00460_));
 sg13g2_inv_1 _07005_ (.Y(_01593_),
    .A(_00332_));
 sg13g2_inv_1 _07006_ (.Y(_01594_),
    .A(_00524_));
 sg13g2_inv_1 _07007_ (.Y(_01595_),
    .A(_00172_));
 sg13g2_inv_1 _07008_ (.Y(_01596_),
    .A(_00461_));
 sg13g2_inv_1 _07009_ (.Y(_01597_),
    .A(_00173_));
 sg13g2_inv_1 _07010_ (.Y(_01598_),
    .A(_00301_));
 sg13g2_inv_1 _07011_ (.Y(_01599_),
    .A(_00206_));
 sg13g2_inv_1 _07012_ (.Y(_01600_),
    .A(_00462_));
 sg13g2_inv_1 _07013_ (.Y(_01601_),
    .A(_00334_));
 sg13g2_inv_1 _07014_ (.Y(_01602_),
    .A(_00430_));
 sg13g2_inv_1 _07015_ (.Y(_01603_),
    .A(_00174_));
 sg13g2_inv_1 _07016_ (.Y(_01604_),
    .A(_00302_));
 sg13g2_inv_1 _07017_ (.Y(_01605_),
    .A(_00207_));
 sg13g2_inv_1 _07018_ (.Y(_01606_),
    .A(_00463_));
 sg13g2_inv_1 _07019_ (.Y(_01607_),
    .A(_00335_));
 sg13g2_inv_1 _07020_ (.Y(_01608_),
    .A(_00175_));
 sg13g2_inv_1 _07021_ (.Y(_01609_),
    .A(_00303_));
 sg13g2_inv_1 _07022_ (.Y(_01610_),
    .A(_00208_));
 sg13g2_inv_1 _07023_ (.Y(_01611_),
    .A(_00464_));
 sg13g2_inv_1 _07024_ (.Y(_01612_),
    .A(_00336_));
 sg13g2_inv_1 _07025_ (.Y(_01613_),
    .A(_00432_));
 sg13g2_inv_1 _07026_ (.Y(_01614_),
    .A(_00176_));
 sg13g2_inv_1 _07027_ (.Y(_01615_),
    .A(_00304_));
 sg13g2_inv_1 _07028_ (.Y(_01616_),
    .A(_00209_));
 sg13g2_inv_1 _07029_ (.Y(_01617_),
    .A(_00465_));
 sg13g2_inv_1 _07030_ (.Y(_01618_),
    .A(_00337_));
 sg13g2_inv_1 _07031_ (.Y(_01619_),
    .A(_00433_));
 sg13g2_inv_1 _07032_ (.Y(_01620_),
    .A(_00177_));
 sg13g2_inv_1 _07033_ (.Y(_01621_),
    .A(_00305_));
 sg13g2_inv_1 _07034_ (.Y(_01622_),
    .A(_00210_));
 sg13g2_inv_1 _07035_ (.Y(_01623_),
    .A(_00466_));
 sg13g2_inv_1 _07036_ (.Y(_01624_),
    .A(_00338_));
 sg13g2_inv_1 _07037_ (.Y(_01625_),
    .A(_00434_));
 sg13g2_inv_1 _07038_ (.Y(_01626_),
    .A(_00178_));
 sg13g2_inv_1 _07039_ (.Y(_01627_),
    .A(_00306_));
 sg13g2_inv_1 _07040_ (.Y(_01628_),
    .A(_00211_));
 sg13g2_inv_1 _07041_ (.Y(_01629_),
    .A(_00467_));
 sg13g2_inv_1 _07042_ (.Y(_01630_),
    .A(_00339_));
 sg13g2_inv_1 _07043_ (.Y(_01631_),
    .A(_00435_));
 sg13g2_inv_1 _07044_ (.Y(_01632_),
    .A(_00179_));
 sg13g2_inv_1 _07045_ (.Y(_01633_),
    .A(_00307_));
 sg13g2_inv_1 _07046_ (.Y(_01634_),
    .A(_00212_));
 sg13g2_inv_1 _07047_ (.Y(_01635_),
    .A(_00468_));
 sg13g2_inv_1 _07048_ (.Y(_01636_),
    .A(_00340_));
 sg13g2_inv_1 _07049_ (.Y(_01637_),
    .A(_00180_));
 sg13g2_inv_1 _07050_ (.Y(_01638_),
    .A(_00308_));
 sg13g2_inv_1 _07051_ (.Y(_01639_),
    .A(_00213_));
 sg13g2_inv_1 _07052_ (.Y(_01640_),
    .A(_00469_));
 sg13g2_inv_1 _07053_ (.Y(_01641_),
    .A(_00341_));
 sg13g2_inv_1 _07054_ (.Y(_01642_),
    .A(_00437_));
 sg13g2_inv_1 _07055_ (.Y(_01643_),
    .A(_00181_));
 sg13g2_inv_1 _07056_ (.Y(_01644_),
    .A(_00309_));
 sg13g2_inv_1 _07057_ (.Y(_01645_),
    .A(_00214_));
 sg13g2_inv_1 _07058_ (.Y(_01646_),
    .A(_00470_));
 sg13g2_inv_1 _07059_ (.Y(_01647_),
    .A(_00342_));
 sg13g2_inv_1 _07060_ (.Y(_01648_),
    .A(_00438_));
 sg13g2_inv_1 _07061_ (.Y(_01649_),
    .A(_00182_));
 sg13g2_inv_1 _07062_ (.Y(_01650_),
    .A(_00310_));
 sg13g2_inv_1 _07063_ (.Y(_01651_),
    .A(\cpu.Bimm[6] ));
 sg13g2_inv_1 _07064_ (.Y(_01652_),
    .A(_00215_));
 sg13g2_inv_1 _07065_ (.Y(_01653_),
    .A(_00471_));
 sg13g2_inv_1 _07066_ (.Y(_01654_),
    .A(_00343_));
 sg13g2_inv_1 _07067_ (.Y(_01655_),
    .A(_00439_));
 sg13g2_inv_1 _07068_ (.Y(_01656_),
    .A(_00183_));
 sg13g2_inv_1 _07069_ (.Y(_01657_),
    .A(_00311_));
 sg13g2_inv_1 _07070_ (.Y(_01658_),
    .A(_00216_));
 sg13g2_inv_1 _07071_ (.Y(_01659_),
    .A(_00472_));
 sg13g2_inv_1 _07072_ (.Y(_01660_),
    .A(_00344_));
 sg13g2_inv_1 _07073_ (.Y(_01661_),
    .A(_00440_));
 sg13g2_inv_1 _07074_ (.Y(_01662_),
    .A(_00184_));
 sg13g2_inv_1 _07075_ (.Y(_01663_),
    .A(_00312_));
 sg13g2_inv_1 _07076_ (.Y(_01664_),
    .A(_00557_));
 sg13g2_inv_1 _07077_ (.Y(_01665_),
    .A(_00217_));
 sg13g2_inv_1 _07078_ (.Y(_01666_),
    .A(_00473_));
 sg13g2_inv_1 _07079_ (.Y(_01667_),
    .A(_00345_));
 sg13g2_inv_1 _07080_ (.Y(_01668_),
    .A(_00441_));
 sg13g2_inv_1 _07081_ (.Y(_01669_),
    .A(_00185_));
 sg13g2_inv_1 _07082_ (.Y(_01670_),
    .A(_00313_));
 sg13g2_inv_1 _07083_ (.Y(_01671_),
    .A(_00218_));
 sg13g2_inv_1 _07084_ (.Y(_01672_),
    .A(_00474_));
 sg13g2_inv_1 _07085_ (.Y(_01673_),
    .A(_00346_));
 sg13g2_inv_1 _07086_ (.Y(_01674_),
    .A(_00442_));
 sg13g2_inv_1 _07087_ (.Y(_01675_),
    .A(_00186_));
 sg13g2_inv_1 _07088_ (.Y(_01676_),
    .A(_00314_));
 sg13g2_inv_1 _07089_ (.Y(_01677_),
    .A(_00219_));
 sg13g2_inv_1 _07090_ (.Y(_01678_),
    .A(_00315_));
 sg13g2_inv_1 _07091_ (.Y(_01679_),
    .A(\cpu.Bimm[2] ));
 sg13g2_inv_1 _07092_ (.Y(_01680_),
    .A(_00156_));
 sg13g2_inv_1 _07093_ (.Y(_01681_),
    .A(_00220_));
 sg13g2_inv_1 _07094_ (.Y(_01682_),
    .A(_00476_));
 sg13g2_inv_1 _07095_ (.Y(_01683_),
    .A(_00348_));
 sg13g2_inv_1 _07096_ (.Y(_01684_),
    .A(_00444_));
 sg13g2_inv_1 _07097_ (.Y(_01685_),
    .A(_00188_));
 sg13g2_inv_1 _07098_ (.Y(_01686_),
    .A(_00316_));
 sg13g2_inv_1 _07099_ (.Y(_01687_),
    .A(\cpu.regs[12][0] ));
 sg13g2_inv_1 _07100_ (.Y(_01688_),
    .A(\cpu.regs[14][0] ));
 sg13g2_inv_1 _07101_ (.Y(_01689_),
    .A(_00189_));
 sg13g2_inv_2 _07102_ (.Y(_01690_),
    .A(\cpu.Bimm[11] ));
 sg13g2_inv_1 _07103_ (.Y(_01691_),
    .A(net3631));
 sg13g2_inv_1 _07104_ (.Y(_01692_),
    .A(_00447_));
 sg13g2_inv_1 _07105_ (.Y(_01693_),
    .A(_00319_));
 sg13g2_inv_1 _07106_ (.Y(_01694_),
    .A(_00415_));
 sg13g2_inv_2 _07107_ (.Y(_01695_),
    .A(net3702));
 sg13g2_inv_1 _07108_ (.Y(_01696_),
    .A(\cpu.IR[4] ));
 sg13g2_inv_4 _07109_ (.A(net3699),
    .Y(_01697_));
 sg13g2_inv_1 _07110_ (.Y(_01698_),
    .A(net3698));
 sg13g2_inv_1 _07111_ (.Y(_01699_),
    .A(\jtag0.tapst[1] ));
 sg13g2_inv_1 _07112_ (.Y(_01700_),
    .A(\jtag0.tapst[3] ));
 sg13g2_inv_1 _07113_ (.Y(_01701_),
    .A(\uart0.txdiv[0] ));
 sg13g2_inv_1 _07114_ (.Y(_01702_),
    .A(\pwmc[1] ));
 sg13g2_inv_1 _07115_ (.Y(_01703_),
    .A(\pwmc[3] ));
 sg13g2_inv_1 _07116_ (.Y(_01704_),
    .A(\pwmc[5] ));
 sg13g2_inv_1 _07117_ (.Y(_01705_),
    .A(_00125_));
 sg13g2_inv_2 _07118_ (.Y(_01706_),
    .A(pwmout));
 sg13g2_inv_1 _07119_ (.Y(_01707_),
    .A(\ckd[0] ));
 sg13g2_inv_1 _07120_ (.Y(_01708_),
    .A(_00197_));
 sg13g2_inv_1 _07121_ (.Y(_01709_),
    .A(_00165_));
 sg13g2_inv_1 _07122_ (.Y(_01710_),
    .A(_00196_));
 sg13g2_inv_1 _07123_ (.Y(_01711_),
    .A(_00452_));
 sg13g2_inv_1 _07124_ (.Y(_01712_),
    .A(_00324_));
 sg13g2_inv_1 _07125_ (.Y(_01713_),
    .A(_00420_));
 sg13g2_inv_1 _07126_ (.Y(_01714_),
    .A(_00164_));
 sg13g2_inv_1 _07127_ (.Y(_01715_),
    .A(_00065_));
 sg13g2_inv_1 _07128_ (.Y(_01716_),
    .A(_00195_));
 sg13g2_inv_1 _07129_ (.Y(_01717_),
    .A(_00163_));
 sg13g2_inv_1 _07130_ (.Y(_01718_),
    .A(_00064_));
 sg13g2_inv_1 _07131_ (.Y(_01719_),
    .A(_00194_));
 sg13g2_inv_1 _07132_ (.Y(_01720_),
    .A(_00199_));
 sg13g2_inv_1 _07133_ (.Y(_01721_),
    .A(_00423_));
 sg13g2_inv_1 _07134_ (.Y(_01722_),
    .A(_00198_));
 sg13g2_inv_1 _07135_ (.Y(_01723_),
    .A(_00422_));
 sg13g2_inv_1 _07136_ (.Y(_01724_),
    .A(_00166_));
 sg13g2_inv_2 _07137_ (.Y(_01725_),
    .A(_00563_));
 sg13g2_inv_1 _07138_ (.Y(_01726_),
    .A(_00564_));
 sg13g2_inv_1 _07139_ (.Y(_01727_),
    .A(_00568_));
 sg13g2_inv_1 _07140_ (.Y(_01728_),
    .A(_00569_));
 sg13g2_inv_4 _07141_ (.A(net3686),
    .Y(_01729_));
 sg13g2_inv_2 _07142_ (.Y(_01730_),
    .A(net3674));
 sg13g2_inv_1 _07143_ (.Y(_01731_),
    .A(\cpu.PCci[17] ));
 sg13g2_inv_1 _07144_ (.Y(_01732_),
    .A(net3655));
 sg13g2_inv_1 _07145_ (.Y(_01733_),
    .A(\irqvect[3][25] ));
 sg13g2_inv_1 _07146_ (.Y(_01734_),
    .A(net914));
 sg13g2_inv_1 _07147_ (.Y(_01735_),
    .A(\tcount[3] ));
 sg13g2_inv_1 _07148_ (.Y(_01736_),
    .A(\tcount[19] ));
 sg13g2_inv_1 _07149_ (.Y(_01737_),
    .A(\tcount[7] ));
 sg13g2_inv_1 _07150_ (.Y(_01738_),
    .A(\tcount[25] ));
 sg13g2_inv_1 _07151_ (.Y(_01739_),
    .A(\tcount[10] ));
 sg13g2_inv_1 _07152_ (.Y(_01740_),
    .A(\tcount[13] ));
 sg13g2_inv_1 _07153_ (.Y(_01741_),
    .A(\uart0.txsh[2] ));
 sg13g2_inv_1 _07154_ (.Y(_01742_),
    .A(\uart0.txsh[3] ));
 sg13g2_inv_1 _07155_ (.Y(_01743_),
    .A(\uart0.txsh[4] ));
 sg13g2_inv_1 _07156_ (.Y(_01744_),
    .A(\uart0.txsh[5] ));
 sg13g2_inv_1 _07157_ (.Y(_01745_),
    .A(\uart0.txsh[6] ));
 sg13g2_inv_1 _07158_ (.Y(_01746_),
    .A(\uart0.txsh[7] ));
 sg13g2_inv_1 _07159_ (.Y(_01747_),
    .A(\uart0.txsh[8] ));
 sg13g2_inv_1 _07160_ (.Y(_01748_),
    .A(\jtag0.stms ));
 sg13g2_inv_1 _07161_ (.Y(_01749_),
    .A(_00124_));
 sg13g2_inv_1 _07162_ (.Y(_00591_),
    .A(net3941));
 sg13g2_nand2b_2 _07163_ (.Y(_01750_),
    .B(\jtag0.tapst[3] ),
    .A_N(net3926));
 sg13g2_nor2_1 _07164_ (.A(_01699_),
    .B(_01750_),
    .Y(_01751_));
 sg13g2_nand2_1 _07165_ (.Y(_01752_),
    .A(net3927),
    .B(\jtag0.tapst[1] ));
 sg13g2_nor2_2 _07166_ (.A(_01750_),
    .B(_01752_),
    .Y(_01753_));
 sg13g2_mux2_1 _07167_ (.A0(\jtag0.irsh[2] ),
    .A1(\jtag0.stdi ),
    .S(_01753_),
    .X(_01534_));
 sg13g2_mux2_1 _07168_ (.A0(\jtag0.irsh[1] ),
    .A1(\jtag0.irsh[2] ),
    .S(_01753_),
    .X(_01533_));
 sg13g2_nand2_1 _07169_ (.Y(_01754_),
    .A(\jtag0.irsh[1] ),
    .B(_01753_));
 sg13g2_o21ai_1 _07170_ (.B1(_01754_),
    .Y(_01532_),
    .A1(_01539_),
    .A2(_01753_));
 sg13g2_nand3b_1 _07171_ (.B(\cpu.IR[1] ),
    .C(\cpu.IR[0] ),
    .Y(_01755_),
    .A_N(\cpu.IR[2] ));
 sg13g2_or2_1 _07172_ (.X(_01756_),
    .B(_00546_),
    .A(\cpu.IR[3] ));
 sg13g2_nand2b_1 _07173_ (.Y(_01757_),
    .B(\cpu.IR[5] ),
    .A_N(\cpu.IR[4] ));
 sg13g2_nor4_2 _07174_ (.A(\cpu.IR[6] ),
    .B(_01755_),
    .C(_01756_),
    .Y(_01758_),
    .D(_01757_));
 sg13g2_nand2b_2 _07175_ (.Y(_01759_),
    .B(net3704),
    .A_N(\cpu.IR[3] ));
 sg13g2_or2_1 _07176_ (.X(_01760_),
    .B(_01759_),
    .A(_01755_));
 sg13g2_or2_1 _07177_ (.X(_01761_),
    .B(\cpu.IR[5] ),
    .A(\cpu.IR[6] ));
 sg13g2_nor3_2 _07178_ (.A(_01755_),
    .B(_01759_),
    .C(_01761_),
    .Y(_01762_));
 sg13g2_nor4_1 _07179_ (.A(\cpu.IR[4] ),
    .B(_01755_),
    .C(_01759_),
    .D(_01761_),
    .Y(_01763_));
 sg13g2_nand2_2 _07180_ (.Y(_01764_),
    .A(_01696_),
    .B(_01762_));
 sg13g2_nor2_1 _07181_ (.A(_01758_),
    .B(net3448),
    .Y(_01765_));
 sg13g2_or2_1 _07182_ (.X(_01766_),
    .B(net3448),
    .A(_01758_));
 sg13g2_mux2_2 _07183_ (.A0(\cpu.PCreg0[31] ),
    .A1(\cpu.PCreg1[31] ),
    .S(net3631),
    .X(\cpu.PC[31] ));
 sg13g2_and2_1 _07184_ (.A(net3406),
    .B(\cpu.PC[31] ),
    .X(_01767_));
 sg13g2_and2_1 _07185_ (.A(net3702),
    .B(net3683),
    .X(_01768_));
 sg13g2_nand2_2 _07186_ (.Y(_01769_),
    .A(net3703),
    .B(net3681));
 sg13g2_mux4_1 _07187_ (.S0(net3577),
    .A0(_00127_),
    .A1(_00191_),
    .A2(_00511_),
    .A3(_00415_),
    .S1(net3655),
    .X(_01770_));
 sg13g2_nor2_1 _07188_ (.A(net3660),
    .B(_01770_),
    .Y(_01771_));
 sg13g2_and2_2 _07189_ (.A(net3704),
    .B(\cpu.IR[18] ),
    .X(_01772_));
 sg13g2_nand2_1 _07190_ (.Y(_01773_),
    .A(net3704),
    .B(\cpu.IR[18] ));
 sg13g2_a221oi_1 _07191_ (.B2(_01693_),
    .C1(net3655),
    .B1(net3588),
    .A1(_01692_),
    .Y(_01774_),
    .A2(net3680));
 sg13g2_nor2_1 _07192_ (.A(_00287_),
    .B(net3618),
    .Y(_01775_));
 sg13g2_o21ai_1 _07193_ (.B1(net3657),
    .Y(_01776_),
    .A1(_00159_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07194_ (.B1(net3669),
    .Y(_01777_),
    .A1(_01775_),
    .A2(_01776_));
 sg13g2_o21ai_1 _07195_ (.B1(net3573),
    .Y(_01778_),
    .A1(_01774_),
    .A2(_01777_));
 sg13g2_nor2_1 _07196_ (.A(_01771_),
    .B(_01778_),
    .Y(_01779_));
 sg13g2_nor2_1 _07197_ (.A(_01695_),
    .B(net3622),
    .Y(_01780_));
 sg13g2_nand2_2 _07198_ (.Y(_01781_),
    .A(net3700),
    .B(net3654));
 sg13g2_nor2_2 _07199_ (.A(\cpu.IR[18] ),
    .B(net3569),
    .Y(_01782_));
 sg13g2_nor2_1 _07200_ (.A(_01695_),
    .B(_01730_),
    .Y(_01783_));
 sg13g2_nand2_1 _07201_ (.Y(_01784_),
    .A(net3703),
    .B(net3665));
 sg13g2_mux4_1 _07202_ (.S0(net3574),
    .A0(_00383_),
    .A1(_00255_),
    .A2(_00223_),
    .A3(_00093_),
    .S1(net3554),
    .X(_01785_));
 sg13g2_nor2_2 _07203_ (.A(net3573),
    .B(net3446),
    .Y(_01786_));
 sg13g2_o21ai_1 _07204_ (.B1(net3554),
    .Y(_01787_),
    .A1(_00479_),
    .A2(net3574));
 sg13g2_nor2_1 _07205_ (.A(_00351_),
    .B(net3680),
    .Y(_01788_));
 sg13g2_a21oi_1 _07206_ (.A1(_00061_),
    .A2(net3662),
    .Y(_01789_),
    .B1(net3574));
 sg13g2_o21ai_1 _07207_ (.B1(_01787_),
    .Y(_01790_),
    .A1(_01788_),
    .A2(_01789_));
 sg13g2_a221oi_1 _07208_ (.B2(_01790_),
    .C1(_01779_),
    .B1(net3396),
    .A1(net3441),
    .Y(_01791_),
    .A2(_01785_));
 sg13g2_nand2_1 _07209_ (.Y(_01792_),
    .A(net3641),
    .B(_01791_));
 sg13g2_a21oi_1 _07210_ (.A1(_01602_),
    .A2(net3598),
    .Y(_01793_),
    .B1(net3670));
 sg13g2_o21ai_1 _07211_ (.B1(_01793_),
    .Y(_01794_),
    .A1(_00526_),
    .A2(net3598));
 sg13g2_a22oi_1 _07212_ (.Y(_01795_),
    .B1(net3598),
    .B2(_01604_),
    .A2(net3690),
    .A1(_01603_));
 sg13g2_a21oi_1 _07213_ (.A1(net3670),
    .A2(_01795_),
    .Y(_01796_),
    .B1(net3620));
 sg13g2_a21oi_1 _07214_ (.A1(_01599_),
    .A2(net3598),
    .Y(_01797_),
    .B1(net3670));
 sg13g2_o21ai_1 _07215_ (.B1(_01797_),
    .Y(_01798_),
    .A1(_00142_),
    .A2(net3598));
 sg13g2_a22oi_1 _07216_ (.Y(_01799_),
    .B1(net3598),
    .B2(_01601_),
    .A2(net3690),
    .A1(_01600_));
 sg13g2_a21oi_1 _07217_ (.A1(net3670),
    .A2(_01799_),
    .Y(_01800_),
    .B1(net3656));
 sg13g2_a221oi_1 _07218_ (.B2(_01800_),
    .C1(net3570),
    .B1(_01798_),
    .A1(_01794_),
    .Y(_01801_),
    .A2(_01796_));
 sg13g2_mux4_1 _07219_ (.S0(net3600),
    .A0(_00398_),
    .A1(_00270_),
    .A2(_00238_),
    .A3(_00108_),
    .S1(net3564),
    .X(_01802_));
 sg13g2_o21ai_1 _07220_ (.B1(net3564),
    .Y(_01803_),
    .A1(_00494_),
    .A2(net3600));
 sg13g2_nor2_1 _07221_ (.A(_00366_),
    .B(net3690),
    .Y(_01804_));
 sg13g2_a21oi_1 _07222_ (.A1(_00076_),
    .A2(net3670),
    .Y(_01805_),
    .B1(net3600));
 sg13g2_o21ai_1 _07223_ (.B1(_01803_),
    .Y(_01806_),
    .A1(_01804_),
    .A2(_01805_));
 sg13g2_a221oi_1 _07224_ (.B2(net3399),
    .C1(_01801_),
    .B1(_01806_),
    .A1(net3444),
    .Y(_01807_),
    .A2(_01802_));
 sg13g2_nor2_2 _07225_ (.A(net3642),
    .B(_01807_),
    .Y(_01808_));
 sg13g2_and2_1 _07226_ (.A(net3642),
    .B(_01807_),
    .X(_01809_));
 sg13g2_a21oi_1 _07227_ (.A1(_01605_),
    .A2(net3599),
    .Y(_01810_),
    .B1(net3670));
 sg13g2_o21ai_1 _07228_ (.B1(_01810_),
    .Y(_01811_),
    .A1(_00143_),
    .A2(net3599));
 sg13g2_a22oi_1 _07229_ (.Y(_01812_),
    .B1(net3599),
    .B2(_01607_),
    .A2(net3690),
    .A1(_01606_));
 sg13g2_a21oi_1 _07230_ (.A1(net3673),
    .A2(_01812_),
    .Y(_01813_),
    .B1(net3656));
 sg13g2_mux2_1 _07231_ (.A0(_00527_),
    .A1(_00431_),
    .S(net3599),
    .X(_01814_));
 sg13g2_a22oi_1 _07232_ (.Y(_01815_),
    .B1(net3599),
    .B2(_01609_),
    .A2(net3690),
    .A1(_01608_));
 sg13g2_nand2_1 _07233_ (.Y(_01816_),
    .A(net3673),
    .B(_01815_));
 sg13g2_a21oi_1 _07234_ (.A1(net3623),
    .A2(_01814_),
    .Y(_01817_),
    .B1(net3620));
 sg13g2_a221oi_1 _07235_ (.B2(_01817_),
    .C1(net3570),
    .B1(_01816_),
    .A1(_01811_),
    .Y(_01818_),
    .A2(_01813_));
 sg13g2_mux4_1 _07236_ (.S0(net3600),
    .A0(_00399_),
    .A1(_00271_),
    .A2(_00239_),
    .A3(_00109_),
    .S1(net3564),
    .X(_01819_));
 sg13g2_o21ai_1 _07237_ (.B1(net3564),
    .Y(_01820_),
    .A1(_00495_),
    .A2(net3598));
 sg13g2_nor2_1 _07238_ (.A(_00367_),
    .B(net3690),
    .Y(_01821_));
 sg13g2_a21oi_1 _07239_ (.A1(_00077_),
    .A2(net3670),
    .Y(_01822_),
    .B1(net3598));
 sg13g2_o21ai_1 _07240_ (.B1(_01820_),
    .Y(_01823_),
    .A1(_01821_),
    .A2(_01822_));
 sg13g2_a221oi_1 _07241_ (.B2(net3399),
    .C1(_01818_),
    .B1(_01823_),
    .A1(net3444),
    .Y(_01824_),
    .A2(_01819_));
 sg13g2_a21oi_1 _07242_ (.A1(_01625_),
    .A2(net3607),
    .Y(_01825_),
    .B1(net3674));
 sg13g2_o21ai_1 _07243_ (.B1(_01825_),
    .Y(_01826_),
    .A1(_00530_),
    .A2(net3607));
 sg13g2_a22oi_1 _07244_ (.Y(_01827_),
    .B1(net3607),
    .B2(_01627_),
    .A2(net3691),
    .A1(_01626_));
 sg13g2_a21oi_1 _07245_ (.A1(net3674),
    .A2(_01827_),
    .Y(_01828_),
    .B1(net3620));
 sg13g2_a21oi_1 _07246_ (.A1(_01622_),
    .A2(net3607),
    .Y(_01829_),
    .B1(net3674));
 sg13g2_o21ai_1 _07247_ (.B1(_01829_),
    .Y(_01830_),
    .A1(_00146_),
    .A2(net3607));
 sg13g2_a22oi_1 _07248_ (.Y(_01831_),
    .B1(net3607),
    .B2(_01624_),
    .A2(net3691),
    .A1(_01623_));
 sg13g2_a21oi_1 _07249_ (.A1(net3674),
    .A2(_01831_),
    .Y(_01832_),
    .B1(net3658));
 sg13g2_a221oi_1 _07250_ (.B2(_01832_),
    .C1(net3570),
    .B1(_01830_),
    .A1(_01826_),
    .Y(_01833_),
    .A2(_01828_));
 sg13g2_mux4_1 _07251_ (.S0(net3608),
    .A0(_00402_),
    .A1(_00274_),
    .A2(_00242_),
    .A3(_00112_),
    .S1(net3567),
    .X(_01834_));
 sg13g2_o21ai_1 _07252_ (.B1(net3566),
    .Y(_01835_),
    .A1(_00498_),
    .A2(net3608));
 sg13g2_nor2_1 _07253_ (.A(_00370_),
    .B(net3691),
    .Y(_01836_));
 sg13g2_a21oi_1 _07254_ (.A1(_00080_),
    .A2(net3674),
    .Y(_01837_),
    .B1(net3607));
 sg13g2_o21ai_1 _07255_ (.B1(_01835_),
    .Y(_01838_),
    .A1(_01836_),
    .A2(_01837_));
 sg13g2_a221oi_1 _07256_ (.B2(net3400),
    .C1(_01833_),
    .B1(_01838_),
    .A1(net3445),
    .Y(_01839_),
    .A2(_01834_));
 sg13g2_xnor2_1 _07257_ (.Y(_01840_),
    .A(net3643),
    .B(_01839_));
 sg13g2_a21oi_1 _07258_ (.A1(_01645_),
    .A2(net3609),
    .Y(_01841_),
    .B1(net3671));
 sg13g2_o21ai_1 _07259_ (.B1(_01841_),
    .Y(_01842_),
    .A1(_00150_),
    .A2(net3609));
 sg13g2_a22oi_1 _07260_ (.Y(_01843_),
    .B1(net3609),
    .B2(_01647_),
    .A2(net3689),
    .A1(_01646_));
 sg13g2_a21oi_1 _07261_ (.A1(net3671),
    .A2(_01843_),
    .Y(_01844_),
    .B1(net3656));
 sg13g2_a21oi_1 _07262_ (.A1(_01648_),
    .A2(net3609),
    .Y(_01845_),
    .B1(net3672));
 sg13g2_o21ai_1 _07263_ (.B1(_01845_),
    .Y(_01846_),
    .A1(_00534_),
    .A2(net3609));
 sg13g2_a22oi_1 _07264_ (.Y(_01847_),
    .B1(net3609),
    .B2(_01650_),
    .A2(net3689),
    .A1(_01649_));
 sg13g2_a21oi_1 _07265_ (.A1(net3671),
    .A2(_01847_),
    .Y(_01848_),
    .B1(net3620));
 sg13g2_a221oi_1 _07266_ (.B2(_01848_),
    .C1(net3570),
    .B1(_01846_),
    .A1(_01842_),
    .Y(_01849_),
    .A2(_01844_));
 sg13g2_mux4_1 _07267_ (.S0(net3602),
    .A0(_00406_),
    .A1(_00278_),
    .A2(_00246_),
    .A3(_00116_),
    .S1(net3565),
    .X(_01850_));
 sg13g2_o21ai_1 _07268_ (.B1(net3565),
    .Y(_01851_),
    .A1(_00502_),
    .A2(net3602));
 sg13g2_nor2_1 _07269_ (.A(_00374_),
    .B(net3689),
    .Y(_01852_));
 sg13g2_a21oi_1 _07270_ (.A1(_00084_),
    .A2(net3672),
    .Y(_01853_),
    .B1(net3602));
 sg13g2_o21ai_1 _07271_ (.B1(_01851_),
    .Y(_01854_),
    .A1(_01852_),
    .A2(_01853_));
 sg13g2_a221oi_1 _07272_ (.B2(net3399),
    .C1(_01849_),
    .B1(_01854_),
    .A1(net3444),
    .Y(_01855_),
    .A2(_01850_));
 sg13g2_nand2b_1 _07273_ (.Y(_01856_),
    .B(_01855_),
    .A_N(_00559_));
 sg13g2_a21oi_1 _07274_ (.A1(_01658_),
    .A2(net3610),
    .Y(_01857_),
    .B1(net3676));
 sg13g2_o21ai_1 _07275_ (.B1(_01857_),
    .Y(_01858_),
    .A1(_00152_),
    .A2(net3610));
 sg13g2_a22oi_1 _07276_ (.Y(_01859_),
    .B1(net3610),
    .B2(_01660_),
    .A2(net3691),
    .A1(_01659_));
 sg13g2_a21oi_1 _07277_ (.A1(net3676),
    .A2(_01859_),
    .Y(_01860_),
    .B1(net3656));
 sg13g2_a21oi_1 _07278_ (.A1(_01661_),
    .A2(net3609),
    .Y(_01861_),
    .B1(net3676));
 sg13g2_o21ai_1 _07279_ (.B1(_01861_),
    .Y(_01862_),
    .A1(_00536_),
    .A2(net3609));
 sg13g2_a22oi_1 _07280_ (.Y(_01863_),
    .B1(net3610),
    .B2(_01663_),
    .A2(net3691),
    .A1(_01662_));
 sg13g2_a21oi_1 _07281_ (.A1(net3676),
    .A2(_01863_),
    .Y(_01864_),
    .B1(net3620));
 sg13g2_a221oi_1 _07282_ (.B2(_01864_),
    .C1(net3570),
    .B1(_01862_),
    .A1(_01858_),
    .Y(_01865_),
    .A2(_01860_));
 sg13g2_mux4_1 _07283_ (.S0(net3603),
    .A0(_00408_),
    .A1(_00280_),
    .A2(_00248_),
    .A3(_00118_),
    .S1(net3565),
    .X(_01866_));
 sg13g2_o21ai_1 _07284_ (.B1(net3565),
    .Y(_01867_),
    .A1(_00504_),
    .A2(net3604));
 sg13g2_nor2_1 _07285_ (.A(_00376_),
    .B(net3689),
    .Y(_01868_));
 sg13g2_a21oi_1 _07286_ (.A1(_00086_),
    .A2(net3672),
    .Y(_01869_),
    .B1(net3604));
 sg13g2_o21ai_1 _07287_ (.B1(_01867_),
    .Y(_01870_),
    .A1(_01868_),
    .A2(_01869_));
 sg13g2_a221oi_1 _07288_ (.B2(net3399),
    .C1(_01865_),
    .B1(_01870_),
    .A1(net3444),
    .Y(_01871_),
    .A2(_01866_));
 sg13g2_nor2_1 _07289_ (.A(_01664_),
    .B(_01871_),
    .Y(_01872_));
 sg13g2_a21oi_1 _07290_ (.A1(_01665_),
    .A2(net3582),
    .Y(_01873_),
    .B1(net3665));
 sg13g2_o21ai_1 _07291_ (.B1(_01873_),
    .Y(_01874_),
    .A1(_00153_),
    .A2(net3578));
 sg13g2_a22oi_1 _07292_ (.Y(_01875_),
    .B1(net3580),
    .B2(_01667_),
    .A2(net3681),
    .A1(_01666_));
 sg13g2_a21oi_1 _07293_ (.A1(net3665),
    .A2(_01875_),
    .Y(_01876_),
    .B1(net3654));
 sg13g2_a21oi_1 _07294_ (.A1(_01668_),
    .A2(net3578),
    .Y(_01877_),
    .B1(net3665));
 sg13g2_o21ai_1 _07295_ (.B1(_01877_),
    .Y(_01878_),
    .A1(_00537_),
    .A2(net3578));
 sg13g2_a22oi_1 _07296_ (.Y(_01879_),
    .B1(net3580),
    .B2(_01670_),
    .A2(net3681),
    .A1(_01669_));
 sg13g2_a21oi_1 _07297_ (.A1(net3665),
    .A2(_01879_),
    .Y(_01880_),
    .B1(net3621));
 sg13g2_a221oi_1 _07298_ (.B2(_01880_),
    .C1(net3571),
    .B1(_01878_),
    .A1(_01874_),
    .Y(_01881_),
    .A2(_01876_));
 sg13g2_mux4_1 _07299_ (.S0(net3579),
    .A0(_00409_),
    .A1(_00281_),
    .A2(_00249_),
    .A3(_00119_),
    .S1(net3556),
    .X(_01882_));
 sg13g2_o21ai_1 _07300_ (.B1(net3556),
    .Y(_01883_),
    .A1(_00505_),
    .A2(net3579));
 sg13g2_nor2_1 _07301_ (.A(_00377_),
    .B(net3681),
    .Y(_01884_));
 sg13g2_a21oi_1 _07302_ (.A1(_00087_),
    .A2(net3665),
    .Y(_01885_),
    .B1(net3579));
 sg13g2_o21ai_1 _07303_ (.B1(_01883_),
    .Y(_01886_),
    .A1(_01884_),
    .A2(_01885_));
 sg13g2_a221oi_1 _07304_ (.B2(net3397),
    .C1(_01881_),
    .B1(_01886_),
    .A1(net3441),
    .Y(_01887_),
    .A2(_01882_));
 sg13g2_inv_1 _07305_ (.Y(_01888_),
    .A(_01887_));
 sg13g2_mux2_1 _07306_ (.A0(_00551_),
    .A1(_00556_),
    .S(net3449),
    .X(_01889_));
 sg13g2_nor2_1 _07307_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sg13g2_a21oi_1 _07308_ (.A1(_01671_),
    .A2(net3603),
    .Y(_01891_),
    .B1(net3671));
 sg13g2_o21ai_1 _07309_ (.B1(_01891_),
    .Y(_01892_),
    .A1(_00154_),
    .A2(net3603));
 sg13g2_a22oi_1 _07310_ (.Y(_01893_),
    .B1(net3603),
    .B2(_01673_),
    .A2(net3693),
    .A1(_01672_));
 sg13g2_a21oi_1 _07311_ (.A1(net3671),
    .A2(_01893_),
    .Y(_01894_),
    .B1(net3656));
 sg13g2_a21oi_1 _07312_ (.A1(_01674_),
    .A2(net3603),
    .Y(_01895_),
    .B1(net3671));
 sg13g2_o21ai_1 _07313_ (.B1(_01895_),
    .Y(_01896_),
    .A1(_00538_),
    .A2(net3603));
 sg13g2_a22oi_1 _07314_ (.Y(_01897_),
    .B1(net3603),
    .B2(_01676_),
    .A2(net3693),
    .A1(_01675_));
 sg13g2_a21oi_1 _07315_ (.A1(net3671),
    .A2(_01897_),
    .Y(_01898_),
    .B1(net3620));
 sg13g2_a221oi_1 _07316_ (.B2(_01898_),
    .C1(net3571),
    .B1(_01896_),
    .A1(_01892_),
    .Y(_01899_),
    .A2(_01894_));
 sg13g2_mux4_1 _07317_ (.S0(net3581),
    .A0(_00410_),
    .A1(_00282_),
    .A2(_00250_),
    .A3(_00120_),
    .S1(net3565),
    .X(_01900_));
 sg13g2_o21ai_1 _07318_ (.B1(net3565),
    .Y(_01901_),
    .A1(_00506_),
    .A2(net3601));
 sg13g2_nor2_1 _07319_ (.A(_00378_),
    .B(net3689),
    .Y(_01902_));
 sg13g2_a21oi_1 _07320_ (.A1(_00088_),
    .A2(net3672),
    .Y(_01903_),
    .B1(net3601));
 sg13g2_o21ai_1 _07321_ (.B1(_01901_),
    .Y(_01904_),
    .A1(_01902_),
    .A2(_01903_));
 sg13g2_a221oi_1 _07322_ (.B2(net3399),
    .C1(_01899_),
    .B1(_01904_),
    .A1(net3444),
    .Y(_01905_),
    .A2(_01900_));
 sg13g2_mux2_1 _07323_ (.A0(_00550_),
    .A1(_00555_),
    .S(net3449),
    .X(_01906_));
 sg13g2_inv_1 _07324_ (.Y(_01907_),
    .A(_01906_));
 sg13g2_nand2_1 _07325_ (.Y(_01908_),
    .A(_01905_),
    .B(_01907_));
 sg13g2_mux2_1 _07326_ (.A0(_00539_),
    .A1(_00443_),
    .S(net3579),
    .X(_01909_));
 sg13g2_nand2b_1 _07327_ (.Y(_01910_),
    .B(net3684),
    .A_N(_00187_));
 sg13g2_a21oi_1 _07328_ (.A1(_01678_),
    .A2(net3578),
    .Y(_01911_),
    .B1(net3556));
 sg13g2_a221oi_1 _07329_ (.B2(_01911_),
    .C1(_01781_),
    .B1(_01910_),
    .A1(net3556),
    .Y(_01912_),
    .A2(_01909_));
 sg13g2_mux2_1 _07330_ (.A0(_00155_),
    .A1(_00219_),
    .S(net3578),
    .X(_01913_));
 sg13g2_a21oi_1 _07331_ (.A1(net3700),
    .A2(net3684),
    .Y(_01914_),
    .B1(_00347_));
 sg13g2_nor2b_1 _07332_ (.A(_00475_),
    .B_N(net3681),
    .Y(_01915_));
 sg13g2_nor3_1 _07333_ (.A(net3556),
    .B(_01914_),
    .C(_01915_),
    .Y(_01916_));
 sg13g2_a221oi_1 _07334_ (.B2(_01913_),
    .C1(_01916_),
    .B1(net3556),
    .A1(net3700),
    .Y(_01917_),
    .A2(net3654));
 sg13g2_or3_1 _07335_ (.A(net3571),
    .B(_01912_),
    .C(_01917_),
    .X(_01918_));
 sg13g2_mux4_1 _07336_ (.S0(net3579),
    .A0(_00411_),
    .A1(_00283_),
    .A2(_00251_),
    .A3(_00121_),
    .S1(net3556),
    .X(_01919_));
 sg13g2_nand2_1 _07337_ (.Y(_01920_),
    .A(net3441),
    .B(_01919_));
 sg13g2_o21ai_1 _07338_ (.B1(net3558),
    .Y(_01921_),
    .A1(_00507_),
    .A2(net3578));
 sg13g2_nor2_1 _07339_ (.A(_00379_),
    .B(net3681),
    .Y(_01922_));
 sg13g2_a21oi_1 _07340_ (.A1(_00089_),
    .A2(net3665),
    .Y(_01923_),
    .B1(net3578));
 sg13g2_o21ai_1 _07341_ (.B1(_01921_),
    .Y(_01924_),
    .A1(_01922_),
    .A2(_01923_));
 sg13g2_nand2_1 _07342_ (.Y(_01925_),
    .A(net3396),
    .B(_01924_));
 sg13g2_and3_2 _07343_ (.X(_01926_),
    .A(_01918_),
    .B(_01920_),
    .C(_01925_));
 sg13g2_nand3_1 _07344_ (.B(_01920_),
    .C(_01925_),
    .A(_01918_),
    .Y(_01927_));
 sg13g2_mux2_1 _07345_ (.A0(_00549_),
    .A1(_00554_),
    .S(net3449),
    .X(_01928_));
 sg13g2_nor2_1 _07346_ (.A(_01927_),
    .B(_01928_),
    .Y(_01929_));
 sg13g2_nand2_1 _07347_ (.Y(_01930_),
    .A(_01927_),
    .B(_01928_));
 sg13g2_nand2b_1 _07348_ (.Y(_01931_),
    .B(_01930_),
    .A_N(_01929_));
 sg13g2_a22oi_1 _07349_ (.Y(_01932_),
    .B1(net3581),
    .B2(_01683_),
    .A2(net3682),
    .A1(_01682_));
 sg13g2_nand2_1 _07350_ (.Y(_01933_),
    .A(_01681_),
    .B(net3581));
 sg13g2_a21oi_1 _07351_ (.A1(_01680_),
    .A2(net3619),
    .Y(_01934_),
    .B1(net3663));
 sg13g2_a221oi_1 _07352_ (.B2(_01934_),
    .C1(net3654),
    .B1(_01933_),
    .A1(net3663),
    .Y(_01935_),
    .A2(_01932_));
 sg13g2_nand2b_1 _07353_ (.Y(_01936_),
    .B(net3619),
    .A_N(_00540_));
 sg13g2_a21oi_1 _07354_ (.A1(_01684_),
    .A2(net3581),
    .Y(_01937_),
    .B1(net3663));
 sg13g2_a22oi_1 _07355_ (.Y(_01938_),
    .B1(net3581),
    .B2(_01686_),
    .A2(net3682),
    .A1(_01685_));
 sg13g2_a221oi_1 _07356_ (.B2(net3663),
    .C1(net3621),
    .B1(_01938_),
    .A1(_01936_),
    .Y(_01939_),
    .A2(_01937_));
 sg13g2_or3_2 _07357_ (.A(net3571),
    .B(_01935_),
    .C(_01939_),
    .X(_01940_));
 sg13g2_mux4_1 _07358_ (.S0(net3580),
    .A0(_00412_),
    .A1(_00284_),
    .A2(_00252_),
    .A3(_00122_),
    .S1(net3557),
    .X(_01941_));
 sg13g2_o21ai_1 _07359_ (.B1(net3557),
    .Y(_01942_),
    .A1(_00508_),
    .A2(net3580));
 sg13g2_nor2_1 _07360_ (.A(_00380_),
    .B(net3682),
    .Y(_01943_));
 sg13g2_a21oi_1 _07361_ (.A1(_00090_),
    .A2(net3663),
    .Y(_01944_),
    .B1(net3580));
 sg13g2_o21ai_1 _07362_ (.B1(_01942_),
    .Y(_01945_),
    .A1(_01943_),
    .A2(_01944_));
 sg13g2_a22oi_1 _07363_ (.Y(_01946_),
    .B1(_01945_),
    .B2(net3397),
    .A2(_01941_),
    .A1(net3442));
 sg13g2_and2_1 _07364_ (.A(_01940_),
    .B(_01946_),
    .X(_01947_));
 sg13g2_or2_1 _07365_ (.X(_01948_),
    .B(net3449),
    .A(_00548_));
 sg13g2_o21ai_1 _07366_ (.B1(_01948_),
    .Y(_01949_),
    .A1(_00553_),
    .A2(_01764_));
 sg13g2_nand3_1 _07367_ (.B(_01946_),
    .C(_01949_),
    .A(_01940_),
    .Y(_01950_));
 sg13g2_mux2_1 _07368_ (.A0(_00157_),
    .A1(_00221_),
    .S(net3580),
    .X(_01951_));
 sg13g2_a21oi_1 _07369_ (.A1(net3702),
    .A2(net3682),
    .Y(_01952_),
    .B1(_00349_));
 sg13g2_nor2b_1 _07370_ (.A(_00477_),
    .B_N(net3682),
    .Y(_01953_));
 sg13g2_nor3_1 _07371_ (.A(net3557),
    .B(_01952_),
    .C(_01953_),
    .Y(_01954_));
 sg13g2_a221oi_1 _07372_ (.B2(_01951_),
    .C1(_01954_),
    .B1(net3557),
    .A1(net3702),
    .Y(_01955_),
    .A2(net3654));
 sg13g2_mux2_1 _07373_ (.A0(_00541_),
    .A1(_00445_),
    .S(net3580),
    .X(_01956_));
 sg13g2_nand2b_1 _07374_ (.Y(_01957_),
    .B(net3580),
    .A_N(_00317_));
 sg13g2_a21oi_1 _07375_ (.A1(_01689_),
    .A2(net3681),
    .Y(_01958_),
    .B1(net3557));
 sg13g2_a221oi_1 _07376_ (.B2(_01958_),
    .C1(_01781_),
    .B1(_01957_),
    .A1(net3557),
    .Y(_01959_),
    .A2(_01956_));
 sg13g2_or3_1 _07377_ (.A(net3571),
    .B(_01955_),
    .C(_01959_),
    .X(_01960_));
 sg13g2_mux4_1 _07378_ (.S0(net3578),
    .A0(_00413_),
    .A1(_00285_),
    .A2(_00253_),
    .A3(_00123_),
    .S1(net3558),
    .X(_01961_));
 sg13g2_nand2_1 _07379_ (.Y(_01962_),
    .A(net3442),
    .B(_01961_));
 sg13g2_o21ai_1 _07380_ (.B1(net3556),
    .Y(_01963_),
    .A1(_00509_),
    .A2(net3579));
 sg13g2_nor2_1 _07381_ (.A(_00381_),
    .B(net3681),
    .Y(_01964_));
 sg13g2_a21oi_1 _07382_ (.A1(_00091_),
    .A2(net3665),
    .Y(_01965_),
    .B1(net3579));
 sg13g2_o21ai_1 _07383_ (.B1(_01963_),
    .Y(_01966_),
    .A1(_01964_),
    .A2(_01965_));
 sg13g2_nand2_1 _07384_ (.Y(_01967_),
    .A(net3396),
    .B(_01966_));
 sg13g2_and3_1 _07385_ (.X(_01968_),
    .A(_01960_),
    .B(_01962_),
    .C(_01967_));
 sg13g2_nand2_1 _07386_ (.Y(_01969_),
    .A(net3645),
    .B(net3449));
 sg13g2_o21ai_1 _07387_ (.B1(_01969_),
    .Y(_01970_),
    .A1(_01690_),
    .A2(net3449));
 sg13g2_nand4_1 _07388_ (.B(_01962_),
    .C(_01967_),
    .A(_01960_),
    .Y(_01971_),
    .D(_01970_));
 sg13g2_a21oi_1 _07389_ (.A1(_01940_),
    .A2(_01946_),
    .Y(_01972_),
    .B1(_01949_));
 sg13g2_o21ai_1 _07390_ (.B1(_01950_),
    .Y(_01973_),
    .A1(_01971_),
    .A2(_01972_));
 sg13g2_a21oi_2 _07391_ (.B1(_01929_),
    .Y(_01974_),
    .A2(_01973_),
    .A1(_01930_));
 sg13g2_xnor2_1 _07392_ (.Y(_01975_),
    .A(_01905_),
    .B(_01907_));
 sg13g2_o21ai_1 _07393_ (.B1(_01908_),
    .Y(_01976_),
    .A1(_01974_),
    .A2(_01975_));
 sg13g2_xnor2_1 _07394_ (.Y(_01977_),
    .A(_01887_),
    .B(_01889_));
 sg13g2_a21oi_1 _07395_ (.A1(_01976_),
    .A2(_01977_),
    .Y(_01978_),
    .B1(_01890_));
 sg13g2_a221oi_1 _07396_ (.B2(_01977_),
    .C1(_01890_),
    .B1(_01976_),
    .A1(_01664_),
    .Y(_01979_),
    .A2(_01871_));
 sg13g2_a21oi_1 _07397_ (.A1(_01655_),
    .A2(net3602),
    .Y(_01980_),
    .B1(net3664));
 sg13g2_o21ai_1 _07398_ (.B1(_01980_),
    .Y(_01981_),
    .A1(_00535_),
    .A2(net3601));
 sg13g2_a22oi_1 _07399_ (.Y(_01982_),
    .B1(net3602),
    .B2(_01657_),
    .A2(net3682),
    .A1(_01656_));
 sg13g2_a21oi_1 _07400_ (.A1(net3663),
    .A2(_01982_),
    .Y(_01983_),
    .B1(net3621));
 sg13g2_a21oi_1 _07401_ (.A1(_01652_),
    .A2(net3601),
    .Y(_01984_),
    .B1(net3664));
 sg13g2_o21ai_1 _07402_ (.B1(_01984_),
    .Y(_01985_),
    .A1(_00151_),
    .A2(net3601));
 sg13g2_a22oi_1 _07403_ (.Y(_01986_),
    .B1(net3581),
    .B2(_01654_),
    .A2(net3682),
    .A1(_01653_));
 sg13g2_a21oi_1 _07404_ (.A1(net3663),
    .A2(_01986_),
    .Y(_01987_),
    .B1(net3654));
 sg13g2_a221oi_1 _07405_ (.B2(_01987_),
    .C1(net3571),
    .B1(_01985_),
    .A1(_01981_),
    .Y(_01988_),
    .A2(_01983_));
 sg13g2_mux4_1 _07406_ (.S0(net3582),
    .A0(_00407_),
    .A1(_00279_),
    .A2(_00247_),
    .A3(_00117_),
    .S1(net3558),
    .X(_01989_));
 sg13g2_o21ai_1 _07407_ (.B1(net3557),
    .Y(_01990_),
    .A1(_00503_),
    .A2(net3582));
 sg13g2_nor2_1 _07408_ (.A(_00375_),
    .B(net3682),
    .Y(_01991_));
 sg13g2_a21oi_1 _07409_ (.A1(_00085_),
    .A2(net3663),
    .Y(_01992_),
    .B1(net3582));
 sg13g2_o21ai_1 _07410_ (.B1(_01990_),
    .Y(_01993_),
    .A1(_01991_),
    .A2(_01992_));
 sg13g2_a221oi_1 _07411_ (.B2(net3397),
    .C1(_01988_),
    .B1(_01993_),
    .A1(net3442),
    .Y(_01994_),
    .A2(_01989_));
 sg13g2_xnor2_1 _07412_ (.Y(_01995_),
    .A(\cpu.Bimm[6] ),
    .B(_01994_));
 sg13g2_nor3_2 _07413_ (.A(_01872_),
    .B(_01979_),
    .C(_01995_),
    .Y(_01996_));
 sg13g2_nor2b_1 _07414_ (.A(_00558_),
    .B_N(_01994_),
    .Y(_01997_));
 sg13g2_xnor2_1 _07415_ (.Y(_01998_),
    .A(_00559_),
    .B(_01855_));
 sg13g2_o21ai_1 _07416_ (.B1(_01998_),
    .Y(_01999_),
    .A1(_01996_),
    .A2(_01997_));
 sg13g2_a21oi_1 _07417_ (.A1(_01639_),
    .A2(net3613),
    .Y(_02000_),
    .B1(net3677));
 sg13g2_o21ai_1 _07418_ (.B1(_02000_),
    .Y(_02001_),
    .A1(_00149_),
    .A2(net3613));
 sg13g2_a22oi_1 _07419_ (.Y(_02002_),
    .B1(net3613),
    .B2(_01641_),
    .A2(net3692),
    .A1(_01640_));
 sg13g2_a21oi_1 _07420_ (.A1(net3677),
    .A2(_02002_),
    .Y(_02003_),
    .B1(net3656));
 sg13g2_a21oi_1 _07421_ (.A1(_01642_),
    .A2(net3612),
    .Y(_02004_),
    .B1(net3677));
 sg13g2_o21ai_1 _07422_ (.B1(_02004_),
    .Y(_02005_),
    .A1(_00533_),
    .A2(net3612));
 sg13g2_a22oi_1 _07423_ (.Y(_02006_),
    .B1(net3611),
    .B2(_01644_),
    .A2(net3692),
    .A1(_01643_));
 sg13g2_a21oi_1 _07424_ (.A1(net3677),
    .A2(_02006_),
    .Y(_02007_),
    .B1(net3620));
 sg13g2_a221oi_1 _07425_ (.B2(_02007_),
    .C1(net3570),
    .B1(_02005_),
    .A1(_02001_),
    .Y(_02008_),
    .A2(_02003_));
 sg13g2_mux4_1 _07426_ (.S0(net3604),
    .A0(_00405_),
    .A1(_00277_),
    .A2(_00245_),
    .A3(_00115_),
    .S1(net3564),
    .X(_02009_));
 sg13g2_o21ai_1 _07427_ (.B1(net3564),
    .Y(_02010_),
    .A1(_00501_),
    .A2(net3604));
 sg13g2_nor2_1 _07428_ (.A(_00373_),
    .B(net3689),
    .Y(_02011_));
 sg13g2_a21oi_1 _07429_ (.A1(_00083_),
    .A2(net3671),
    .Y(_02012_),
    .B1(net3604));
 sg13g2_o21ai_1 _07430_ (.B1(_02010_),
    .Y(_02013_),
    .A1(_02011_),
    .A2(_02012_));
 sg13g2_a221oi_1 _07431_ (.B2(net3399),
    .C1(_02008_),
    .B1(_02013_),
    .A1(net3444),
    .Y(_02014_),
    .A2(_02009_));
 sg13g2_xnor2_1 _07432_ (.Y(_02015_),
    .A(\cpu.Bimm[8] ),
    .B(_02014_));
 sg13g2_a21oi_1 _07433_ (.A1(_01856_),
    .A2(_01999_),
    .Y(_02016_),
    .B1(_02015_));
 sg13g2_nor2b_1 _07434_ (.A(_00560_),
    .B_N(_02014_),
    .Y(_02017_));
 sg13g2_nor2_1 _07435_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sg13g2_a21oi_1 _07436_ (.A1(_01634_),
    .A2(net3601),
    .Y(_02019_),
    .B1(net3672));
 sg13g2_o21ai_1 _07437_ (.B1(_02019_),
    .Y(_02020_),
    .A1(_00148_),
    .A2(net3601));
 sg13g2_a22oi_1 _07438_ (.Y(_02021_),
    .B1(net3601),
    .B2(_01636_),
    .A2(net3689),
    .A1(_01635_));
 sg13g2_a21oi_1 _07439_ (.A1(net3672),
    .A2(_02021_),
    .Y(_02022_),
    .B1(net3656));
 sg13g2_mux2_1 _07440_ (.A0(_00532_),
    .A1(_00436_),
    .S(net3599),
    .X(_02023_));
 sg13g2_a22oi_1 _07441_ (.Y(_02024_),
    .B1(net3603),
    .B2(_01638_),
    .A2(net3689),
    .A1(_01637_));
 sg13g2_nand2_1 _07442_ (.Y(_02025_),
    .A(net3672),
    .B(_02024_));
 sg13g2_a21oi_1 _07443_ (.A1(net3623),
    .A2(_02023_),
    .Y(_02026_),
    .B1(net3621));
 sg13g2_a221oi_1 _07444_ (.B2(_02026_),
    .C1(net3570),
    .B1(_02025_),
    .A1(_02020_),
    .Y(_02027_),
    .A2(_02022_));
 sg13g2_mux4_1 _07445_ (.S0(net3600),
    .A0(_00404_),
    .A1(_00276_),
    .A2(_00244_),
    .A3(_00114_),
    .S1(net3564),
    .X(_02028_));
 sg13g2_o21ai_1 _07446_ (.B1(net3564),
    .Y(_02029_),
    .A1(_00500_),
    .A2(net3600));
 sg13g2_nor2_1 _07447_ (.A(_00372_),
    .B(net3690),
    .Y(_02030_));
 sg13g2_a21oi_1 _07448_ (.A1(_00082_),
    .A2(net3670),
    .Y(_02031_),
    .B1(net3600));
 sg13g2_o21ai_1 _07449_ (.B1(_02029_),
    .Y(_02032_),
    .A1(_02030_),
    .A2(_02031_));
 sg13g2_a221oi_1 _07450_ (.B2(net3399),
    .C1(_02027_),
    .B1(_02032_),
    .A1(net3444),
    .Y(_02033_),
    .A2(_02028_));
 sg13g2_xnor2_1 _07451_ (.Y(_02034_),
    .A(\cpu.Bimm[9] ),
    .B(_02033_));
 sg13g2_inv_1 _07452_ (.Y(_02035_),
    .A(_02034_));
 sg13g2_o21ai_1 _07453_ (.B1(_02035_),
    .Y(_02036_),
    .A1(_02016_),
    .A2(_02017_));
 sg13g2_nand2b_1 _07454_ (.Y(_02037_),
    .B(_02033_),
    .A_N(_00561_));
 sg13g2_and2_1 _07455_ (.A(_02036_),
    .B(_02037_),
    .X(_02038_));
 sg13g2_a21oi_1 _07456_ (.A1(_01631_),
    .A2(net3612),
    .Y(_02039_),
    .B1(net3676));
 sg13g2_o21ai_1 _07457_ (.B1(_02039_),
    .Y(_02040_),
    .A1(_00531_),
    .A2(net3612));
 sg13g2_a22oi_1 _07458_ (.Y(_02041_),
    .B1(net3612),
    .B2(_01633_),
    .A2(net3692),
    .A1(_01632_));
 sg13g2_a21oi_1 _07459_ (.A1(net3676),
    .A2(_02041_),
    .Y(_02042_),
    .B1(net3620));
 sg13g2_a21oi_1 _07460_ (.A1(_01628_),
    .A2(net3612),
    .Y(_02043_),
    .B1(net3677));
 sg13g2_o21ai_1 _07461_ (.B1(_02043_),
    .Y(_02044_),
    .A1(_00147_),
    .A2(net3612));
 sg13g2_a22oi_1 _07462_ (.Y(_02045_),
    .B1(net3612),
    .B2(_01630_),
    .A2(net3692),
    .A1(_01629_));
 sg13g2_a21oi_1 _07463_ (.A1(net3676),
    .A2(_02045_),
    .Y(_02046_),
    .B1(net3656));
 sg13g2_a221oi_1 _07464_ (.B2(_02046_),
    .C1(net3570),
    .B1(_02044_),
    .A1(_02040_),
    .Y(_02047_),
    .A2(_02042_));
 sg13g2_mux4_1 _07465_ (.S0(net3611),
    .A0(_00403_),
    .A1(_00275_),
    .A2(_00243_),
    .A3(_00113_),
    .S1(net3566),
    .X(_02048_));
 sg13g2_o21ai_1 _07466_ (.B1(net3566),
    .Y(_02049_),
    .A1(_00499_),
    .A2(net3611));
 sg13g2_nor2_1 _07467_ (.A(_00371_),
    .B(net3691),
    .Y(_02050_));
 sg13g2_a21oi_1 _07468_ (.A1(_00081_),
    .A2(net3676),
    .Y(_02051_),
    .B1(net3611));
 sg13g2_o21ai_1 _07469_ (.B1(_02049_),
    .Y(_02052_),
    .A1(_02050_),
    .A2(_02051_));
 sg13g2_a221oi_1 _07470_ (.B2(net3399),
    .C1(_02047_),
    .B1(_02052_),
    .A1(net3444),
    .Y(_02053_),
    .A2(_02048_));
 sg13g2_nand2b_1 _07471_ (.Y(_02054_),
    .B(_02053_),
    .A_N(\cpu.Bimm[10] ));
 sg13g2_nand2b_1 _07472_ (.Y(_02055_),
    .B(\cpu.Bimm[10] ),
    .A_N(_02053_));
 sg13g2_and2_1 _07473_ (.A(_02054_),
    .B(_02055_),
    .X(_02056_));
 sg13g2_nor2_1 _07474_ (.A(_02038_),
    .B(_02056_),
    .Y(_02057_));
 sg13g2_nor2b_1 _07475_ (.A(_00562_),
    .B_N(_02053_),
    .Y(_02058_));
 sg13g2_nor2_1 _07476_ (.A(_02057_),
    .B(_02058_),
    .Y(_02059_));
 sg13g2_a221oi_1 _07477_ (.B2(_02055_),
    .C1(_01840_),
    .B1(_02054_),
    .A1(_02036_),
    .Y(_02060_),
    .A2(_02037_));
 sg13g2_nor2b_1 _07478_ (.A(_01840_),
    .B_N(_02058_),
    .Y(_02061_));
 sg13g2_a21o_1 _07479_ (.A2(_01839_),
    .A1(_01575_),
    .B1(_02061_),
    .X(_02062_));
 sg13g2_nor2_1 _07480_ (.A(_02060_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_a21oi_1 _07481_ (.A1(_01619_),
    .A2(net3575),
    .Y(_02064_),
    .B1(net3660));
 sg13g2_o21ai_1 _07482_ (.B1(_02064_),
    .Y(_02065_),
    .A1(_00529_),
    .A2(net3575));
 sg13g2_a22oi_1 _07483_ (.Y(_02066_),
    .B1(net3575),
    .B2(_01621_),
    .A2(net3680),
    .A1(_01620_));
 sg13g2_a21oi_1 _07484_ (.A1(net3661),
    .A2(_02066_),
    .Y(_02067_),
    .B1(net3622));
 sg13g2_a21oi_1 _07485_ (.A1(_01616_),
    .A2(net3577),
    .Y(_02068_),
    .B1(net3660));
 sg13g2_o21ai_1 _07486_ (.B1(_02068_),
    .Y(_02069_),
    .A1(_00145_),
    .A2(net3575));
 sg13g2_a22oi_1 _07487_ (.Y(_02070_),
    .B1(net3576),
    .B2(_01618_),
    .A2(net3685),
    .A1(_01617_));
 sg13g2_a21oi_1 _07488_ (.A1(net3661),
    .A2(_02070_),
    .Y(_02071_),
    .B1(net3655));
 sg13g2_a221oi_1 _07489_ (.B2(_02071_),
    .C1(net3572),
    .B1(_02069_),
    .A1(_02065_),
    .Y(_02072_),
    .A2(_02067_));
 sg13g2_mux4_1 _07490_ (.S0(net3574),
    .A0(_00401_),
    .A1(_00273_),
    .A2(_00241_),
    .A3(_00111_),
    .S1(net3554),
    .X(_02073_));
 sg13g2_o21ai_1 _07491_ (.B1(net3554),
    .Y(_02074_),
    .A1(_00497_),
    .A2(net3576));
 sg13g2_nor2_1 _07492_ (.A(_00369_),
    .B(net3680),
    .Y(_02075_));
 sg13g2_a21oi_1 _07493_ (.A1(_00079_),
    .A2(net3662),
    .Y(_02076_),
    .B1(net3576));
 sg13g2_o21ai_1 _07494_ (.B1(_02074_),
    .Y(_02077_),
    .A1(_02075_),
    .A2(_02076_));
 sg13g2_a221oi_1 _07495_ (.B2(net3396),
    .C1(_02072_),
    .B1(_02077_),
    .A1(net3441),
    .Y(_02078_),
    .A2(_02073_));
 sg13g2_xnor2_1 _07496_ (.Y(_02079_),
    .A(net3643),
    .B(_02078_));
 sg13g2_inv_1 _07497_ (.Y(_02080_),
    .A(_02079_));
 sg13g2_nor2_1 _07498_ (.A(_02063_),
    .B(_02079_),
    .Y(_02081_));
 sg13g2_o21ai_1 _07499_ (.B1(_02080_),
    .Y(_02082_),
    .A1(_02060_),
    .A2(_02062_));
 sg13g2_a21oi_1 _07500_ (.A1(_01610_),
    .A2(net3586),
    .Y(_02083_),
    .B1(net3660));
 sg13g2_o21ai_1 _07501_ (.B1(_02083_),
    .Y(_02084_),
    .A1(_00144_),
    .A2(net3586));
 sg13g2_a22oi_1 _07502_ (.Y(_02085_),
    .B1(net3586),
    .B2(_01612_),
    .A2(net3688),
    .A1(_01611_));
 sg13g2_a21oi_1 _07503_ (.A1(net3669),
    .A2(_02085_),
    .Y(_02086_),
    .B1(net3655));
 sg13g2_a21oi_1 _07504_ (.A1(_01613_),
    .A2(net3585),
    .Y(_02087_),
    .B1(net3660));
 sg13g2_o21ai_1 _07505_ (.B1(_02087_),
    .Y(_02088_),
    .A1(_00528_),
    .A2(net3585));
 sg13g2_a22oi_1 _07506_ (.Y(_02089_),
    .B1(net3585),
    .B2(_01615_),
    .A2(net3688),
    .A1(_01614_));
 sg13g2_a21oi_1 _07507_ (.A1(net3669),
    .A2(_02089_),
    .Y(_02090_),
    .B1(net3622));
 sg13g2_a221oi_1 _07508_ (.B2(_02090_),
    .C1(net3572),
    .B1(_02088_),
    .A1(_02084_),
    .Y(_02091_),
    .A2(_02086_));
 sg13g2_mux4_1 _07509_ (.S0(net3574),
    .A0(_00400_),
    .A1(_00272_),
    .A2(_00240_),
    .A3(_00110_),
    .S1(net3554),
    .X(_02092_));
 sg13g2_o21ai_1 _07510_ (.B1(net3554),
    .Y(_02093_),
    .A1(_00496_),
    .A2(net3574));
 sg13g2_nor2_1 _07511_ (.A(_00368_),
    .B(net3680),
    .Y(_02094_));
 sg13g2_a21oi_1 _07512_ (.A1(_00078_),
    .A2(net3662),
    .Y(_02095_),
    .B1(net3574));
 sg13g2_o21ai_1 _07513_ (.B1(_02093_),
    .Y(_02096_),
    .A1(_02094_),
    .A2(_02095_));
 sg13g2_a221oi_1 _07514_ (.B2(net3396),
    .C1(_02091_),
    .B1(_02096_),
    .A1(net3441),
    .Y(_02097_),
    .A2(_02092_));
 sg13g2_xnor2_1 _07515_ (.Y(_02098_),
    .A(net3642),
    .B(_02097_));
 sg13g2_a21oi_1 _07516_ (.A1(net3642),
    .A2(_02078_),
    .Y(_02099_),
    .B1(_02097_));
 sg13g2_or2_1 _07517_ (.X(_02100_),
    .B(_02099_),
    .A(net3638));
 sg13g2_o21ai_1 _07518_ (.B1(_02100_),
    .Y(_02101_),
    .A1(_02082_),
    .A2(_02098_));
 sg13g2_xnor2_1 _07519_ (.Y(_02102_),
    .A(net3639),
    .B(_01824_));
 sg13g2_a22oi_1 _07520_ (.Y(_02103_),
    .B1(_02101_),
    .B2(_02102_),
    .A2(_01824_),
    .A1(net3642));
 sg13g2_a221oi_1 _07521_ (.B2(_02102_),
    .C1(_01809_),
    .B1(_02101_),
    .A1(net3642),
    .Y(_02104_),
    .A2(_01824_));
 sg13g2_nor2_1 _07522_ (.A(_01808_),
    .B(_01809_),
    .Y(_02105_));
 sg13g2_mux4_1 _07523_ (.S0(net3583),
    .A0(_00141_),
    .A1(_00205_),
    .A2(_00525_),
    .A3(_00429_),
    .S1(net3654),
    .X(_02106_));
 sg13g2_nor2_1 _07524_ (.A(net3664),
    .B(_02106_),
    .Y(_02107_));
 sg13g2_nand2b_1 _07525_ (.Y(_02108_),
    .B(net3600),
    .A_N(_00333_));
 sg13g2_a21oi_1 _07526_ (.A1(_01596_),
    .A2(net3683),
    .Y(_02109_),
    .B1(net3659));
 sg13g2_a22oi_1 _07527_ (.Y(_02110_),
    .B1(net3583),
    .B2(_01598_),
    .A2(net3683),
    .A1(_01597_));
 sg13g2_a221oi_1 _07528_ (.B2(net3654),
    .C1(net3623),
    .B1(_02110_),
    .A1(_02108_),
    .Y(_02111_),
    .A2(_02109_));
 sg13g2_nor3_1 _07529_ (.A(net3571),
    .B(_02107_),
    .C(_02111_),
    .Y(_02112_));
 sg13g2_mux4_1 _07530_ (.S0(net3581),
    .A0(_00397_),
    .A1(_00269_),
    .A2(_00237_),
    .A3(_00107_),
    .S1(net3558),
    .X(_02113_));
 sg13g2_o21ai_1 _07531_ (.B1(net3557),
    .Y(_02114_),
    .A1(_00493_),
    .A2(net3581));
 sg13g2_nor2_1 _07532_ (.A(_00365_),
    .B(net3683),
    .Y(_02115_));
 sg13g2_a21oi_1 _07533_ (.A1(_00075_),
    .A2(net3664),
    .Y(_02116_),
    .B1(net3583));
 sg13g2_o21ai_1 _07534_ (.B1(_02114_),
    .Y(_02117_),
    .A1(_02115_),
    .A2(_02116_));
 sg13g2_a221oi_1 _07535_ (.B2(net3397),
    .C1(_02112_),
    .B1(_02117_),
    .A1(net3442),
    .Y(_02118_),
    .A2(_02113_));
 sg13g2_xnor2_1 _07536_ (.Y(_02119_),
    .A(net3628),
    .B(_02118_));
 sg13g2_nor3_1 _07537_ (.A(_01808_),
    .B(_02104_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_nand2b_1 _07538_ (.Y(_02121_),
    .B(net3616),
    .A_N(_00519_));
 sg13g2_a21oi_1 _07539_ (.A1(_01721_),
    .A2(net3590),
    .Y(_02122_),
    .B1(net3439));
 sg13g2_mux2_1 _07540_ (.A0(_00167_),
    .A1(_00295_),
    .S(net3590),
    .X(_02123_));
 sg13g2_a221oi_1 _07541_ (.B2(net3439),
    .C1(net3569),
    .B1(_02123_),
    .A1(_02121_),
    .Y(_02124_),
    .A2(_02122_));
 sg13g2_mux4_1 _07542_ (.S0(net3590),
    .A0(_00455_),
    .A1(_00327_),
    .A2(_00135_),
    .A3(_00199_),
    .S1(net3562),
    .X(_02125_));
 sg13g2_o21ai_1 _07543_ (.B1(net3573),
    .Y(_02126_),
    .A1(net3446),
    .A2(_02125_));
 sg13g2_mux4_1 _07544_ (.S0(net3593),
    .A0(_00391_),
    .A1(_00263_),
    .A2(_00231_),
    .A3(_00101_),
    .S1(net3563),
    .X(_02127_));
 sg13g2_o21ai_1 _07545_ (.B1(net3563),
    .Y(_02128_),
    .A1(_00487_),
    .A2(net3593));
 sg13g2_nor2_1 _07546_ (.A(_00359_),
    .B(net3686),
    .Y(_02129_));
 sg13g2_a21oi_1 _07547_ (.A1(_00069_),
    .A2(net3667),
    .Y(_02130_),
    .B1(net3593));
 sg13g2_o21ai_1 _07548_ (.B1(_02128_),
    .Y(_02131_),
    .A1(_02129_),
    .A2(_02130_));
 sg13g2_a22oi_1 _07549_ (.Y(_02132_),
    .B1(_02131_),
    .B2(net3400),
    .A2(_02127_),
    .A1(net3445));
 sg13g2_o21ai_1 _07550_ (.B1(_02132_),
    .Y(_02133_),
    .A1(_02124_),
    .A2(_02126_));
 sg13g2_inv_2 _07551_ (.Y(_02134_),
    .A(_02133_));
 sg13g2_xnor2_1 _07552_ (.Y(_02135_),
    .A(net3628),
    .B(_02133_));
 sg13g2_a21oi_1 _07553_ (.A1(_01723_),
    .A2(net3590),
    .Y(_02136_),
    .B1(net3439));
 sg13g2_o21ai_1 _07554_ (.B1(_02136_),
    .Y(_02137_),
    .A1(_00518_),
    .A2(net3590));
 sg13g2_a21oi_1 _07555_ (.A1(_01724_),
    .A2(net3687),
    .Y(_02138_),
    .B1(net3562));
 sg13g2_o21ai_1 _07556_ (.B1(_02138_),
    .Y(_02139_),
    .A1(_00294_),
    .A2(net3616));
 sg13g2_nand3_1 _07557_ (.B(_02137_),
    .C(_02139_),
    .A(net3446),
    .Y(_02140_));
 sg13g2_a21oi_1 _07558_ (.A1(_01722_),
    .A2(net3590),
    .Y(_02141_),
    .B1(net3439));
 sg13g2_o21ai_1 _07559_ (.B1(_02141_),
    .Y(_02142_),
    .A1(_00134_),
    .A2(net3590));
 sg13g2_mux2_1 _07560_ (.A0(_00454_),
    .A1(_00326_),
    .S(net3590),
    .X(_02143_));
 sg13g2_a21oi_1 _07561_ (.A1(net3439),
    .A2(_02143_),
    .Y(_02144_),
    .B1(net3446));
 sg13g2_a21oi_1 _07562_ (.A1(_02142_),
    .A2(_02144_),
    .Y(_02145_),
    .B1(net3572));
 sg13g2_mux4_1 _07563_ (.S0(net3597),
    .A0(_00390_),
    .A1(_00262_),
    .A2(_00230_),
    .A3(_00100_),
    .S1(net3562),
    .X(_02146_));
 sg13g2_and2_1 _07564_ (.A(net3443),
    .B(_02146_),
    .X(_02147_));
 sg13g2_o21ai_1 _07565_ (.B1(net3562),
    .Y(_02148_),
    .A1(_00486_),
    .A2(net3591));
 sg13g2_nor2_1 _07566_ (.A(_00358_),
    .B(net3687),
    .Y(_02149_));
 sg13g2_a21oi_1 _07567_ (.A1(_00068_),
    .A2(net3668),
    .Y(_02150_),
    .B1(net3591));
 sg13g2_o21ai_1 _07568_ (.B1(_02148_),
    .Y(_02151_),
    .A1(_02149_),
    .A2(_02150_));
 sg13g2_a221oi_1 _07569_ (.B2(net3398),
    .C1(_02147_),
    .B1(_02151_),
    .A1(_02140_),
    .Y(_02152_),
    .A2(_02145_));
 sg13g2_xor2_1 _07570_ (.B(_02152_),
    .A(net3643),
    .X(_02153_));
 sg13g2_nand2_1 _07571_ (.Y(_02154_),
    .A(_02135_),
    .B(_02153_));
 sg13g2_o21ai_1 _07572_ (.B1(net3623),
    .Y(_02155_),
    .A1(_00424_),
    .A2(net3616));
 sg13g2_a21oi_1 _07573_ (.A1(_01579_),
    .A2(net3616),
    .Y(_02156_),
    .B1(_02155_));
 sg13g2_nor2_1 _07574_ (.A(_00296_),
    .B(net3616),
    .Y(_02157_));
 sg13g2_o21ai_1 _07575_ (.B1(net3668),
    .Y(_02158_),
    .A1(_00168_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07576_ (.B1(net3657),
    .Y(_02159_),
    .A1(_02157_),
    .A2(_02158_));
 sg13g2_a21oi_1 _07577_ (.A1(_01576_),
    .A2(net3592),
    .Y(_02160_),
    .B1(net3668));
 sg13g2_o21ai_1 _07578_ (.B1(_02160_),
    .Y(_02161_),
    .A1(_00136_),
    .A2(net3592));
 sg13g2_a22oi_1 _07579_ (.Y(_02162_),
    .B1(net3592),
    .B2(_01578_),
    .A2(net3687),
    .A1(_01577_));
 sg13g2_a21oi_1 _07580_ (.A1(net3668),
    .A2(_02162_),
    .Y(_02163_),
    .B1(net3657));
 sg13g2_o21ai_1 _07581_ (.B1(net3573),
    .Y(_02164_),
    .A1(_02156_),
    .A2(_02159_));
 sg13g2_a21oi_1 _07582_ (.A1(_02161_),
    .A2(_02163_),
    .Y(_02165_),
    .B1(_02164_));
 sg13g2_mux4_1 _07583_ (.S0(net3592),
    .A0(_00392_),
    .A1(_00264_),
    .A2(_00232_),
    .A3(_00102_),
    .S1(net3562),
    .X(_02166_));
 sg13g2_o21ai_1 _07584_ (.B1(net3562),
    .Y(_02167_),
    .A1(_00488_),
    .A2(net3597));
 sg13g2_nor2_1 _07585_ (.A(_00360_),
    .B(net3687),
    .Y(_02168_));
 sg13g2_a21oi_1 _07586_ (.A1(_00070_),
    .A2(net3668),
    .Y(_02169_),
    .B1(net3592));
 sg13g2_o21ai_1 _07587_ (.B1(_02167_),
    .Y(_02170_),
    .A1(_02168_),
    .A2(_02169_));
 sg13g2_a221oi_1 _07588_ (.B2(net3398),
    .C1(_02165_),
    .B1(_02170_),
    .A1(net3443),
    .Y(_02171_),
    .A2(_02166_));
 sg13g2_nor2_1 _07589_ (.A(net3638),
    .B(_02171_),
    .Y(_02172_));
 sg13g2_a21oi_1 _07590_ (.A1(_01581_),
    .A2(net3585),
    .Y(_02173_),
    .B1(net3439));
 sg13g2_o21ai_1 _07591_ (.B1(_02173_),
    .Y(_02174_),
    .A1(_00521_),
    .A2(net3585));
 sg13g2_mux2_1 _07592_ (.A0(_00169_),
    .A1(_00297_),
    .S(net3585),
    .X(_02175_));
 sg13g2_a21oi_1 _07593_ (.A1(net3439),
    .A2(_02175_),
    .Y(_02176_),
    .B1(net3569));
 sg13g2_mux4_1 _07594_ (.S0(net3585),
    .A0(_00457_),
    .A1(_00329_),
    .A2(_00137_),
    .A3(_00201_),
    .S1(net3559),
    .X(_02177_));
 sg13g2_o21ai_1 _07595_ (.B1(net3573),
    .Y(_02178_),
    .A1(net3447),
    .A2(_02177_));
 sg13g2_a21oi_1 _07596_ (.A1(_02174_),
    .A2(_02176_),
    .Y(_02179_),
    .B1(_02178_));
 sg13g2_mux4_1 _07597_ (.S0(net3574),
    .A0(_00393_),
    .A1(_00265_),
    .A2(_00233_),
    .A3(_00103_),
    .S1(net3554),
    .X(_02180_));
 sg13g2_o21ai_1 _07598_ (.B1(net3555),
    .Y(_02181_),
    .A1(_00489_),
    .A2(net3576));
 sg13g2_nor2_1 _07599_ (.A(_00361_),
    .B(net3685),
    .Y(_02182_));
 sg13g2_a21oi_1 _07600_ (.A1(_00071_),
    .A2(net3660),
    .Y(_02183_),
    .B1(net3576));
 sg13g2_o21ai_1 _07601_ (.B1(_02181_),
    .Y(_02184_),
    .A1(_02182_),
    .A2(_02183_));
 sg13g2_a221oi_1 _07602_ (.B2(net3396),
    .C1(_02179_),
    .B1(_02184_),
    .A1(net3441),
    .Y(_02185_),
    .A2(_02180_));
 sg13g2_a21oi_1 _07603_ (.A1(net3638),
    .A2(_02185_),
    .Y(_02186_),
    .B1(_02172_));
 sg13g2_nor2b_1 _07604_ (.A(_02171_),
    .B_N(_02185_),
    .Y(_02187_));
 sg13g2_or3_2 _07605_ (.A(_02154_),
    .B(_02186_),
    .C(_02187_),
    .X(_02188_));
 sg13g2_a21oi_1 _07606_ (.A1(_01587_),
    .A2(net3594),
    .Y(_02189_),
    .B1(net3667));
 sg13g2_o21ai_1 _07607_ (.B1(_02189_),
    .Y(_02190_),
    .A1(_00139_),
    .A2(net3594));
 sg13g2_a22oi_1 _07608_ (.Y(_02191_),
    .B1(net3594),
    .B2(_01589_),
    .A2(net3686),
    .A1(_01588_));
 sg13g2_a21oi_1 _07609_ (.A1(net3667),
    .A2(_02191_),
    .Y(_02192_),
    .B1(net3657));
 sg13g2_o21ai_1 _07610_ (.B1(net3623),
    .Y(_02193_),
    .A1(_00523_),
    .A2(net3596));
 sg13g2_a21oi_1 _07611_ (.A1(_01590_),
    .A2(net3596),
    .Y(_02194_),
    .B1(_02193_));
 sg13g2_nor2_1 _07612_ (.A(_00299_),
    .B(net3617),
    .Y(_02195_));
 sg13g2_o21ai_1 _07613_ (.B1(net3666),
    .Y(_02196_),
    .A1(_00171_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07614_ (.B1(net3657),
    .Y(_02197_),
    .A1(_02195_),
    .A2(_02196_));
 sg13g2_o21ai_1 _07615_ (.B1(_01772_),
    .Y(_02198_),
    .A1(_02194_),
    .A2(_02197_));
 sg13g2_a21oi_1 _07616_ (.A1(_02190_),
    .A2(_02192_),
    .Y(_02199_),
    .B1(_02198_));
 sg13g2_mux4_1 _07617_ (.S0(net3594),
    .A0(_00395_),
    .A1(_00267_),
    .A2(_00235_),
    .A3(_00105_),
    .S1(net3561),
    .X(_02200_));
 sg13g2_o21ai_1 _07618_ (.B1(net3561),
    .Y(_02201_),
    .A1(_00491_),
    .A2(net3595));
 sg13g2_nor2_1 _07619_ (.A(_00363_),
    .B(net3686),
    .Y(_02202_));
 sg13g2_a21oi_1 _07620_ (.A1(_00073_),
    .A2(net3666),
    .Y(_02203_),
    .B1(net3594));
 sg13g2_o21ai_1 _07621_ (.B1(_02201_),
    .Y(_02204_),
    .A1(_02202_),
    .A2(_02203_));
 sg13g2_a221oi_1 _07622_ (.B2(net3398),
    .C1(_02199_),
    .B1(_02204_),
    .A1(net3443),
    .Y(_02205_),
    .A2(_02200_));
 sg13g2_o21ai_1 _07623_ (.B1(net3623),
    .Y(_02206_),
    .A1(_00428_),
    .A2(net3619));
 sg13g2_a21oi_1 _07624_ (.A1(_01594_),
    .A2(net3619),
    .Y(_02207_),
    .B1(_02206_));
 sg13g2_nor2_1 _07625_ (.A(_00300_),
    .B(net3619),
    .Y(_02208_));
 sg13g2_o21ai_1 _07626_ (.B1(net3674),
    .Y(_02209_),
    .A1(_00172_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07627_ (.B1(net3658),
    .Y(_02210_),
    .A1(_02208_),
    .A2(_02209_));
 sg13g2_a21oi_1 _07628_ (.A1(_01591_),
    .A2(net3608),
    .Y(_02211_),
    .B1(net3675));
 sg13g2_o21ai_1 _07629_ (.B1(_02211_),
    .Y(_02212_),
    .A1(_00140_),
    .A2(net3614));
 sg13g2_a22oi_1 _07630_ (.Y(_02213_),
    .B1(net3614),
    .B2(_01593_),
    .A2(net3691),
    .A1(_01592_));
 sg13g2_a21oi_1 _07631_ (.A1(net3674),
    .A2(_02213_),
    .Y(_02214_),
    .B1(net3658));
 sg13g2_o21ai_1 _07632_ (.B1(_01772_),
    .Y(_02215_),
    .A1(_02207_),
    .A2(_02210_));
 sg13g2_a21oi_1 _07633_ (.A1(_02212_),
    .A2(_02214_),
    .Y(_02216_),
    .B1(_02215_));
 sg13g2_mux4_1 _07634_ (.S0(net3608),
    .A0(_00396_),
    .A1(_00268_),
    .A2(_00236_),
    .A3(_00106_),
    .S1(net3566),
    .X(_02217_));
 sg13g2_o21ai_1 _07635_ (.B1(net3566),
    .Y(_02218_),
    .A1(_00492_),
    .A2(net3608));
 sg13g2_nor2_1 _07636_ (.A(_00364_),
    .B(net3691),
    .Y(_02219_));
 sg13g2_a21oi_1 _07637_ (.A1(_00074_),
    .A2(net3675),
    .Y(_02220_),
    .B1(net3608));
 sg13g2_o21ai_1 _07638_ (.B1(_02218_),
    .Y(_02221_),
    .A1(_02219_),
    .A2(_02220_));
 sg13g2_a221oi_1 _07639_ (.B2(net3400),
    .C1(_02216_),
    .B1(_02221_),
    .A1(net3445),
    .Y(_02222_),
    .A2(_02217_));
 sg13g2_and2_1 _07640_ (.A(net3639),
    .B(_02222_),
    .X(_02223_));
 sg13g2_nor2_1 _07641_ (.A(net3639),
    .B(_02222_),
    .Y(_02224_));
 sg13g2_mux2_1 _07642_ (.A0(_02224_),
    .A1(_02223_),
    .S(_02205_),
    .X(_02225_));
 sg13g2_o21ai_1 _07643_ (.B1(_01730_),
    .Y(_02226_),
    .A1(_00426_),
    .A2(net3619));
 sg13g2_a21oi_1 _07644_ (.A1(_01585_),
    .A2(net3619),
    .Y(_02227_),
    .B1(_02226_));
 sg13g2_nor2_1 _07645_ (.A(_00298_),
    .B(net3617),
    .Y(_02228_));
 sg13g2_o21ai_1 _07646_ (.B1(net3666),
    .Y(_02229_),
    .A1(_00170_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07647_ (.B1(net3657),
    .Y(_02230_),
    .A1(_02228_),
    .A2(_02229_));
 sg13g2_a21oi_1 _07648_ (.A1(_01582_),
    .A2(net3594),
    .Y(_02231_),
    .B1(net3666));
 sg13g2_o21ai_1 _07649_ (.B1(_02231_),
    .Y(_02232_),
    .A1(_00138_),
    .A2(net3594));
 sg13g2_a22oi_1 _07650_ (.Y(_02233_),
    .B1(net3594),
    .B2(_01584_),
    .A2(net3686),
    .A1(_01583_));
 sg13g2_a21oi_1 _07651_ (.A1(net3666),
    .A2(_02233_),
    .Y(_02234_),
    .B1(net3657));
 sg13g2_o21ai_1 _07652_ (.B1(_01772_),
    .Y(_02235_),
    .A1(_02227_),
    .A2(_02230_));
 sg13g2_a21oi_1 _07653_ (.A1(_02232_),
    .A2(_02234_),
    .Y(_02236_),
    .B1(_02235_));
 sg13g2_mux4_1 _07654_ (.S0(net3593),
    .A0(_00394_),
    .A1(_00266_),
    .A2(_00234_),
    .A3(_00104_),
    .S1(net3561),
    .X(_02237_));
 sg13g2_o21ai_1 _07655_ (.B1(net3566),
    .Y(_02238_),
    .A1(_00490_),
    .A2(net3607));
 sg13g2_nor2_1 _07656_ (.A(_00362_),
    .B(net3686),
    .Y(_02239_));
 sg13g2_a21oi_1 _07657_ (.A1(_00072_),
    .A2(net3675),
    .Y(_02240_),
    .B1(net3608));
 sg13g2_o21ai_1 _07658_ (.B1(_02238_),
    .Y(_02241_),
    .A1(_02239_),
    .A2(_02240_));
 sg13g2_a221oi_1 _07659_ (.B2(net3398),
    .C1(_02236_),
    .B1(_02241_),
    .A1(net3443),
    .Y(_02242_),
    .A2(_02237_));
 sg13g2_xor2_1 _07660_ (.B(_02242_),
    .A(net3642),
    .X(_02243_));
 sg13g2_nand3b_1 _07661_ (.B(_02225_),
    .C(_02243_),
    .Y(_02244_),
    .A_N(_02188_));
 sg13g2_nor4_2 _07662_ (.A(_01808_),
    .B(_02104_),
    .C(_02119_),
    .Y(_02245_),
    .D(_02244_));
 sg13g2_a22oi_1 _07663_ (.Y(_02246_),
    .B1(_02172_),
    .B2(_02185_),
    .A2(_02171_),
    .A1(net3643));
 sg13g2_nor2_1 _07664_ (.A(_02154_),
    .B(_02246_),
    .Y(_02247_));
 sg13g2_nor4_1 _07665_ (.A(_02118_),
    .B(_02205_),
    .C(_02222_),
    .D(_02242_),
    .Y(_02248_));
 sg13g2_nor2_1 _07666_ (.A(_02134_),
    .B(_02152_),
    .Y(_02249_));
 sg13g2_o21ai_1 _07667_ (.B1(_02249_),
    .Y(_02250_),
    .A1(_02188_),
    .A2(_02248_));
 sg13g2_a21o_1 _07668_ (.A2(_02250_),
    .A1(net3643),
    .B1(_02247_),
    .X(_02251_));
 sg13g2_nor2_1 _07669_ (.A(_00514_),
    .B(net3593),
    .Y(_02252_));
 sg13g2_o21ai_1 _07670_ (.B1(net3561),
    .Y(_02253_),
    .A1(_00418_),
    .A2(net3616));
 sg13g2_mux2_1 _07671_ (.A0(_00162_),
    .A1(_00290_),
    .S(net3593),
    .X(_02254_));
 sg13g2_a21oi_1 _07672_ (.A1(net3440),
    .A2(_02254_),
    .Y(_02255_),
    .B1(net3569));
 sg13g2_o21ai_1 _07673_ (.B1(_02255_),
    .Y(_02256_),
    .A1(_02252_),
    .A2(_02253_));
 sg13g2_a21oi_1 _07674_ (.A1(_01719_),
    .A2(net3591),
    .Y(_02257_),
    .B1(net3440));
 sg13g2_o21ai_1 _07675_ (.B1(_02257_),
    .Y(_02258_),
    .A1(_00130_),
    .A2(net3591));
 sg13g2_mux2_1 _07676_ (.A0(_00450_),
    .A1(_00322_),
    .S(net3591),
    .X(_02259_));
 sg13g2_a21oi_1 _07677_ (.A1(net3440),
    .A2(_02259_),
    .Y(_02260_),
    .B1(net3446));
 sg13g2_a21oi_1 _07678_ (.A1(_02258_),
    .A2(_02260_),
    .Y(_02261_),
    .B1(net3572));
 sg13g2_mux4_1 _07679_ (.S0(net3587),
    .A0(_00386_),
    .A1(_00258_),
    .A2(_00226_),
    .A3(_00096_),
    .S1(net3561),
    .X(_02262_));
 sg13g2_and2_1 _07680_ (.A(net3445),
    .B(_02262_),
    .X(_02263_));
 sg13g2_o21ai_1 _07681_ (.B1(net3561),
    .Y(_02264_),
    .A1(_00482_),
    .A2(net3593));
 sg13g2_nor2_1 _07682_ (.A(_00354_),
    .B(net3686),
    .Y(_02265_));
 sg13g2_a21oi_1 _07683_ (.A1(_00064_),
    .A2(net3667),
    .Y(_02266_),
    .B1(net3593));
 sg13g2_o21ai_1 _07684_ (.B1(_02264_),
    .Y(_02267_),
    .A1(_02265_),
    .A2(_02266_));
 sg13g2_a221oi_1 _07685_ (.B2(net3400),
    .C1(_02263_),
    .B1(_02267_),
    .A1(_02256_),
    .Y(_02268_),
    .A2(_02261_));
 sg13g2_xor2_1 _07686_ (.B(_02268_),
    .A(net3641),
    .X(_02269_));
 sg13g2_mux2_1 _07687_ (.A0(_00515_),
    .A1(_00419_),
    .S(net3585),
    .X(_02270_));
 sg13g2_a21oi_1 _07688_ (.A1(_01717_),
    .A2(net3688),
    .Y(_02271_),
    .B1(net3559));
 sg13g2_o21ai_1 _07689_ (.B1(_02271_),
    .Y(_02272_),
    .A1(_00291_),
    .A2(net3618));
 sg13g2_a21oi_1 _07690_ (.A1(net3559),
    .A2(_02270_),
    .Y(_02273_),
    .B1(net3569));
 sg13g2_mux4_1 _07691_ (.S0(net3575),
    .A0(_00451_),
    .A1(_00323_),
    .A2(_00131_),
    .A3(_00195_),
    .S1(net3559),
    .X(_02274_));
 sg13g2_o21ai_1 _07692_ (.B1(net3573),
    .Y(_02275_),
    .A1(net3447),
    .A2(_02274_));
 sg13g2_a21oi_1 _07693_ (.A1(_02272_),
    .A2(_02273_),
    .Y(_02276_),
    .B1(_02275_));
 sg13g2_mux4_1 _07694_ (.S0(net3575),
    .A0(_00387_),
    .A1(_00259_),
    .A2(_00227_),
    .A3(_00097_),
    .S1(net3555),
    .X(_02277_));
 sg13g2_o21ai_1 _07695_ (.B1(net3555),
    .Y(_02278_),
    .A1(_00483_),
    .A2(net3575));
 sg13g2_nor2_1 _07696_ (.A(_00355_),
    .B(net3680),
    .Y(_02279_));
 sg13g2_a21oi_1 _07697_ (.A1(_00065_),
    .A2(net3660),
    .Y(_02280_),
    .B1(net3575));
 sg13g2_o21ai_1 _07698_ (.B1(_02278_),
    .Y(_02281_),
    .A1(_02279_),
    .A2(_02280_));
 sg13g2_a221oi_1 _07699_ (.B2(net3396),
    .C1(_02276_),
    .B1(_02281_),
    .A1(net3441),
    .Y(_02282_),
    .A2(_02277_));
 sg13g2_xnor2_1 _07700_ (.Y(_02283_),
    .A(net3638),
    .B(_02282_));
 sg13g2_nand2_1 _07701_ (.Y(_02284_),
    .A(_02269_),
    .B(_02283_));
 sg13g2_mux2_1 _07702_ (.A0(_00517_),
    .A1(_00421_),
    .S(net3586),
    .X(_02285_));
 sg13g2_a21oi_1 _07703_ (.A1(_01709_),
    .A2(net3688),
    .Y(_02286_),
    .B1(net3559));
 sg13g2_o21ai_1 _07704_ (.B1(_02286_),
    .Y(_02287_),
    .A1(_00293_),
    .A2(net3616));
 sg13g2_a21oi_1 _07705_ (.A1(net3559),
    .A2(_02285_),
    .Y(_02288_),
    .B1(net3569));
 sg13g2_mux4_1 _07706_ (.S0(net3589),
    .A0(_00453_),
    .A1(_00325_),
    .A2(_00133_),
    .A3(_00197_),
    .S1(net3562),
    .X(_02289_));
 sg13g2_o21ai_1 _07707_ (.B1(net3573),
    .Y(_02290_),
    .A1(net3446),
    .A2(_02289_));
 sg13g2_a21oi_1 _07708_ (.A1(_02287_),
    .A2(_02288_),
    .Y(_02291_),
    .B1(_02290_));
 sg13g2_mux4_1 _07709_ (.S0(net3586),
    .A0(_00389_),
    .A1(_00261_),
    .A2(_00229_),
    .A3(_00099_),
    .S1(net3559),
    .X(_02292_));
 sg13g2_o21ai_1 _07710_ (.B1(net3560),
    .Y(_02293_),
    .A1(_00485_),
    .A2(net3587));
 sg13g2_nor2_1 _07711_ (.A(_00357_),
    .B(net3688),
    .Y(_02294_));
 sg13g2_a21oi_1 _07712_ (.A1(_00067_),
    .A2(net3669),
    .Y(_02295_),
    .B1(net3587));
 sg13g2_o21ai_1 _07713_ (.B1(_02293_),
    .Y(_02296_),
    .A1(_02294_),
    .A2(_02295_));
 sg13g2_a221oi_1 _07714_ (.B2(net3398),
    .C1(_02291_),
    .B1(_02296_),
    .A1(net3443),
    .Y(_02297_),
    .A2(_02292_));
 sg13g2_and2_1 _07715_ (.A(net3628),
    .B(_02297_),
    .X(_02298_));
 sg13g2_nor2_1 _07716_ (.A(_00516_),
    .B(net3595),
    .Y(_02299_));
 sg13g2_a21oi_1 _07717_ (.A1(_01713_),
    .A2(net3595),
    .Y(_02300_),
    .B1(_02299_));
 sg13g2_a21oi_1 _07718_ (.A1(_01714_),
    .A2(net3687),
    .Y(_02301_),
    .B1(net3623));
 sg13g2_o21ai_1 _07719_ (.B1(_02301_),
    .Y(_02302_),
    .A1(_00292_),
    .A2(net3617));
 sg13g2_a21oi_1 _07720_ (.A1(net3623),
    .A2(_02300_),
    .Y(_02303_),
    .B1(net3622));
 sg13g2_a21oi_1 _07721_ (.A1(_01710_),
    .A2(net3595),
    .Y(_02304_),
    .B1(net3666));
 sg13g2_o21ai_1 _07722_ (.B1(_02304_),
    .Y(_02305_),
    .A1(_00132_),
    .A2(net3595));
 sg13g2_a22oi_1 _07723_ (.Y(_02306_),
    .B1(net3595),
    .B2(_01712_),
    .A2(net3686),
    .A1(_01711_));
 sg13g2_a21oi_1 _07724_ (.A1(net3666),
    .A2(_02306_),
    .Y(_02307_),
    .B1(net3657));
 sg13g2_a221oi_1 _07725_ (.B2(_02307_),
    .C1(net3572),
    .B1(_02305_),
    .A1(_02302_),
    .Y(_02308_),
    .A2(_02303_));
 sg13g2_mux4_1 _07726_ (.S0(net3592),
    .A0(_00388_),
    .A1(_00260_),
    .A2(_00228_),
    .A3(_00098_),
    .S1(net3562),
    .X(_02309_));
 sg13g2_o21ai_1 _07727_ (.B1(net3563),
    .Y(_02310_),
    .A1(_00484_),
    .A2(net3595));
 sg13g2_nor2_1 _07728_ (.A(_00356_),
    .B(net3687),
    .Y(_02311_));
 sg13g2_a21oi_1 _07729_ (.A1(_00066_),
    .A2(net3666),
    .Y(_02312_),
    .B1(net3595));
 sg13g2_o21ai_1 _07730_ (.B1(_02310_),
    .Y(_02313_),
    .A1(_02311_),
    .A2(_02312_));
 sg13g2_a221oi_1 _07731_ (.B2(net3398),
    .C1(_02308_),
    .B1(_02313_),
    .A1(net3443),
    .Y(_02314_),
    .A2(_02309_));
 sg13g2_nor2_1 _07732_ (.A(net3638),
    .B(_02314_),
    .Y(_02315_));
 sg13g2_a21oi_1 _07733_ (.A1(_02297_),
    .A2(_02314_),
    .Y(_02316_),
    .B1(_02315_));
 sg13g2_nor3_1 _07734_ (.A(_02284_),
    .B(_02298_),
    .C(_02316_),
    .Y(_02317_));
 sg13g2_o21ai_1 _07735_ (.B1(_02317_),
    .Y(_02318_),
    .A1(_02245_),
    .A2(_02251_));
 sg13g2_a21oi_1 _07736_ (.A1(net3641),
    .A2(_02314_),
    .Y(_02319_),
    .B1(_02298_));
 sg13g2_nand3b_1 _07737_ (.B(_02282_),
    .C(net3641),
    .Y(_02320_),
    .A_N(_02268_));
 sg13g2_o21ai_1 _07738_ (.B1(_02320_),
    .Y(_02321_),
    .A1(_02284_),
    .A2(_02319_));
 sg13g2_a21oi_1 _07739_ (.A1(net3628),
    .A2(_02268_),
    .Y(_02322_),
    .B1(_02321_));
 sg13g2_nor2_1 _07740_ (.A(_00513_),
    .B(net3586),
    .Y(_02323_));
 sg13g2_o21ai_1 _07741_ (.B1(net3559),
    .Y(_02324_),
    .A1(_00417_),
    .A2(net3616));
 sg13g2_mux2_1 _07742_ (.A0(_00161_),
    .A1(_00289_),
    .S(net3586),
    .X(_02325_));
 sg13g2_o21ai_1 _07743_ (.B1(net3446),
    .Y(_02326_),
    .A1(_02323_),
    .A2(_02324_));
 sg13g2_a21oi_1 _07744_ (.A1(net3440),
    .A2(_02325_),
    .Y(_02327_),
    .B1(_02326_));
 sg13g2_mux2_1 _07745_ (.A0(_00129_),
    .A1(_00193_),
    .S(net3587),
    .X(_02328_));
 sg13g2_nor2_1 _07746_ (.A(_00321_),
    .B(net3618),
    .Y(_02329_));
 sg13g2_o21ai_1 _07747_ (.B1(net3440),
    .Y(_02330_),
    .A1(_00449_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07748_ (.B1(net3569),
    .Y(_02331_),
    .A1(_02329_),
    .A2(_02330_));
 sg13g2_a21oi_1 _07749_ (.A1(net3560),
    .A2(_02328_),
    .Y(_02332_),
    .B1(_02331_));
 sg13g2_nor3_1 _07750_ (.A(net3572),
    .B(_02327_),
    .C(_02332_),
    .Y(_02333_));
 sg13g2_mux4_1 _07751_ (.S0(net3588),
    .A0(_00385_),
    .A1(_00257_),
    .A2(_00225_),
    .A3(_00095_),
    .S1(net3560),
    .X(_02334_));
 sg13g2_o21ai_1 _07752_ (.B1(net3560),
    .Y(_02335_),
    .A1(_00481_),
    .A2(net3588));
 sg13g2_nor2_1 _07753_ (.A(_00353_),
    .B(net3688),
    .Y(_02336_));
 sg13g2_a21oi_1 _07754_ (.A1(_00063_),
    .A2(net3669),
    .Y(_02337_),
    .B1(net3588));
 sg13g2_o21ai_1 _07755_ (.B1(_02335_),
    .Y(_02338_),
    .A1(_02336_),
    .A2(_02337_));
 sg13g2_a221oi_1 _07756_ (.B2(net3398),
    .C1(_02333_),
    .B1(_02338_),
    .A1(net3443),
    .Y(_02339_),
    .A2(_02334_));
 sg13g2_xnor2_1 _07757_ (.Y(_02340_),
    .A(net3628),
    .B(_02339_));
 sg13g2_a21o_1 _07758_ (.A2(_02322_),
    .A1(_02318_),
    .B1(_02340_),
    .X(_02341_));
 sg13g2_nor2_1 _07759_ (.A(_00512_),
    .B(net3587),
    .Y(_02342_));
 sg13g2_o21ai_1 _07760_ (.B1(net3561),
    .Y(_02343_),
    .A1(_00416_),
    .A2(net3617));
 sg13g2_mux2_1 _07761_ (.A0(_00160_),
    .A1(_00288_),
    .S(net3596),
    .X(_02344_));
 sg13g2_o21ai_1 _07762_ (.B1(net3447),
    .Y(_02345_),
    .A1(_02342_),
    .A2(_02343_));
 sg13g2_a21oi_1 _07763_ (.A1(net3440),
    .A2(_02344_),
    .Y(_02346_),
    .B1(_02345_));
 sg13g2_mux2_1 _07764_ (.A0(_00128_),
    .A1(_00192_),
    .S(net3596),
    .X(_02347_));
 sg13g2_nor2_1 _07765_ (.A(_00320_),
    .B(net3617),
    .Y(_02348_));
 sg13g2_o21ai_1 _07766_ (.B1(net3440),
    .Y(_02349_),
    .A1(_00448_),
    .A2(_01729_));
 sg13g2_o21ai_1 _07767_ (.B1(net3569),
    .Y(_02350_),
    .A1(_02348_),
    .A2(_02349_));
 sg13g2_a21oi_1 _07768_ (.A1(net3561),
    .A2(_02347_),
    .Y(_02351_),
    .B1(_02350_));
 sg13g2_nor3_1 _07769_ (.A(net3572),
    .B(_02346_),
    .C(_02351_),
    .Y(_02352_));
 sg13g2_mux4_1 _07770_ (.S0(net3587),
    .A0(_00384_),
    .A1(_00256_),
    .A2(_00224_),
    .A3(_00094_),
    .S1(net3560),
    .X(_02353_));
 sg13g2_o21ai_1 _07771_ (.B1(net3560),
    .Y(_02354_),
    .A1(_00480_),
    .A2(net3587));
 sg13g2_nor2_1 _07772_ (.A(_00352_),
    .B(net3688),
    .Y(_02355_));
 sg13g2_a21oi_1 _07773_ (.A1(_00062_),
    .A2(net3669),
    .Y(_02356_),
    .B1(net3587));
 sg13g2_o21ai_1 _07774_ (.B1(_02354_),
    .Y(_02357_),
    .A1(_02355_),
    .A2(_02356_));
 sg13g2_a221oi_1 _07775_ (.B2(net3398),
    .C1(_02352_),
    .B1(_02357_),
    .A1(net3443),
    .Y(_02358_),
    .A2(_02353_));
 sg13g2_nand2_1 _07776_ (.Y(_02359_),
    .A(net3638),
    .B(_02358_));
 sg13g2_or2_1 _07777_ (.X(_02360_),
    .B(_02358_),
    .A(net3638));
 sg13g2_nand2_1 _07778_ (.Y(_02361_),
    .A(_02359_),
    .B(_02360_));
 sg13g2_inv_1 _07779_ (.Y(_02362_),
    .A(_02361_));
 sg13g2_a221oi_1 _07780_ (.B2(_02360_),
    .C1(_02340_),
    .B1(_02359_),
    .A1(_02318_),
    .Y(_02363_),
    .A2(_02322_));
 sg13g2_a21oi_1 _07781_ (.A1(net3628),
    .A2(_02339_),
    .Y(_02364_),
    .B1(_02358_));
 sg13g2_nand2b_1 _07782_ (.Y(_02365_),
    .B(net3641),
    .A_N(_02364_));
 sg13g2_inv_1 _07783_ (.Y(_02366_),
    .A(_02365_));
 sg13g2_xor2_1 _07784_ (.B(_01791_),
    .A(net3641),
    .X(_02367_));
 sg13g2_o21ai_1 _07785_ (.B1(_02367_),
    .Y(_02368_),
    .A1(_02363_),
    .A2(_02366_));
 sg13g2_nor2_1 _07786_ (.A(_00510_),
    .B(net3589),
    .Y(_02369_));
 sg13g2_o21ai_1 _07787_ (.B1(net3560),
    .Y(_02370_),
    .A1(_00414_),
    .A2(net3618));
 sg13g2_mux2_1 _07788_ (.A0(_00158_),
    .A1(_00286_),
    .S(net3589),
    .X(_02371_));
 sg13g2_o21ai_1 _07789_ (.B1(net3446),
    .Y(_02372_),
    .A1(_02369_),
    .A2(_02370_));
 sg13g2_a21oi_2 _07790_ (.B1(_02372_),
    .Y(_02373_),
    .A2(_02371_),
    .A1(net3439));
 sg13g2_mux4_1 _07791_ (.S0(net3577),
    .A0(_00446_),
    .A1(_00318_),
    .A2(_00126_),
    .A3(_00190_),
    .S1(net3555),
    .X(_02374_));
 sg13g2_o21ai_1 _07792_ (.B1(net3573),
    .Y(_02375_),
    .A1(net3447),
    .A2(_02374_));
 sg13g2_mux4_1 _07793_ (.S0(net3584),
    .A0(_00382_),
    .A1(_00254_),
    .A2(_00222_),
    .A3(_00092_),
    .S1(net3554),
    .X(_02376_));
 sg13g2_o21ai_1 _07794_ (.B1(net3555),
    .Y(_02377_),
    .A1(_00478_),
    .A2(net3576));
 sg13g2_nor2_1 _07795_ (.A(_00350_),
    .B(net3685),
    .Y(_02378_));
 sg13g2_a21oi_1 _07796_ (.A1(_00060_),
    .A2(net3660),
    .Y(_02379_),
    .B1(net3576));
 sg13g2_o21ai_1 _07797_ (.B1(_02377_),
    .Y(_02380_),
    .A1(_02378_),
    .A2(_02379_));
 sg13g2_a22oi_1 _07798_ (.Y(_02381_),
    .B1(_02380_),
    .B2(net3396),
    .A2(_02376_),
    .A1(net3441));
 sg13g2_o21ai_1 _07799_ (.B1(_02381_),
    .Y(_02382_),
    .A1(_02373_),
    .A2(_02375_));
 sg13g2_inv_1 _07800_ (.Y(_02383_),
    .A(_02382_));
 sg13g2_xor2_1 _07801_ (.B(_02382_),
    .A(net3641),
    .X(_02384_));
 sg13g2_nand3_1 _07802_ (.B(_02368_),
    .C(_02384_),
    .A(_01792_),
    .Y(_02385_));
 sg13g2_a21o_2 _07803_ (.A2(_02368_),
    .A1(_01792_),
    .B1(_02384_),
    .X(_02386_));
 sg13g2_and3_2 _07804_ (.X(_02387_),
    .A(net3403),
    .B(_02385_),
    .C(_02386_));
 sg13g2_nor2_1 _07805_ (.A(net3405),
    .B(\cpu.PC[31] ),
    .Y(_02388_));
 sg13g2_a21oi_2 _07806_ (.B1(net3407),
    .Y(_02389_),
    .A2(_02386_),
    .A1(_02385_));
 sg13g2_mux2_2 _07807_ (.A0(\cpu.PCreg0[29] ),
    .A1(\cpu.PCreg1[29] ),
    .S(net3631),
    .X(\cpu.PC[29] ));
 sg13g2_nand2_1 _07808_ (.Y(_02390_),
    .A(net3407),
    .B(\cpu.PC[29] ));
 sg13g2_and2_1 _07809_ (.A(net3641),
    .B(_02339_),
    .X(_02391_));
 sg13g2_inv_1 _07810_ (.Y(_02392_),
    .A(_02391_));
 sg13g2_nand3_1 _07811_ (.B(_02362_),
    .C(_02392_),
    .A(_02341_),
    .Y(_02393_));
 sg13g2_a21o_1 _07812_ (.A2(_02392_),
    .A1(_02341_),
    .B1(_02362_),
    .X(_02394_));
 sg13g2_nand3_1 _07813_ (.B(_02393_),
    .C(_02394_),
    .A(net3404),
    .Y(_02395_));
 sg13g2_or2_1 _07814_ (.X(_02396_),
    .B(\cpu.PC[29] ),
    .A(net3404));
 sg13g2_a21o_1 _07815_ (.A2(_02394_),
    .A1(_02393_),
    .B1(net3407),
    .X(_02397_));
 sg13g2_mux2_2 _07816_ (.A0(\cpu.PCreg0[30] ),
    .A1(\cpu.PCreg1[30] ),
    .S(net3631),
    .X(\cpu.PC[30] ));
 sg13g2_nand2_1 _07817_ (.Y(_02398_),
    .A(net3407),
    .B(\cpu.PC[30] ));
 sg13g2_or3_1 _07818_ (.A(_02363_),
    .B(_02366_),
    .C(_02367_),
    .X(_02399_));
 sg13g2_nand3_1 _07819_ (.B(_02368_),
    .C(_02399_),
    .A(net3404),
    .Y(_02400_));
 sg13g2_or2_1 _07820_ (.X(_02401_),
    .B(\cpu.PC[30] ),
    .A(net3404));
 sg13g2_a21o_1 _07821_ (.A2(_02399_),
    .A1(_02368_),
    .B1(net3407),
    .X(_02402_));
 sg13g2_nand4_1 _07822_ (.B(_02397_),
    .C(_02401_),
    .A(_02396_),
    .Y(_02403_),
    .D(_02402_));
 sg13g2_nor3_2 _07823_ (.A(_02388_),
    .B(_02389_),
    .C(_02403_),
    .Y(_02404_));
 sg13g2_mux2_2 _07824_ (.A0(\cpu.PCreg0[7] ),
    .A1(\cpu.PCreg1[7] ),
    .S(net3636),
    .X(\cpu.PC[7] ));
 sg13g2_nand2_1 _07825_ (.Y(_02405_),
    .A(net3407),
    .B(\cpu.PC[7] ));
 sg13g2_nor3_1 _07826_ (.A(_01996_),
    .B(_01997_),
    .C(_01998_),
    .Y(_02406_));
 sg13g2_nand2_1 _07827_ (.Y(_02407_),
    .A(net3405),
    .B(_01999_));
 sg13g2_o21ai_1 _07828_ (.B1(_02405_),
    .Y(_02408_),
    .A1(_02406_),
    .A2(_02407_));
 sg13g2_mux2_2 _07829_ (.A0(\cpu.PCreg0[6] ),
    .A1(\cpu.PCreg1[6] ),
    .S(net3636),
    .X(\cpu.PC[6] ));
 sg13g2_and2_1 _07830_ (.A(net3406),
    .B(\cpu.PC[6] ),
    .X(_02409_));
 sg13g2_o21ai_1 _07831_ (.B1(_01995_),
    .Y(_02410_),
    .A1(_01872_),
    .A2(_01979_));
 sg13g2_nor2_1 _07832_ (.A(net3406),
    .B(_01996_),
    .Y(_02411_));
 sg13g2_a21o_1 _07833_ (.A2(_02411_),
    .A1(_02410_),
    .B1(_02409_),
    .X(_02412_));
 sg13g2_inv_1 _07834_ (.Y(_02413_),
    .A(net3122));
 sg13g2_nand2b_1 _07835_ (.Y(_02414_),
    .B(net3118),
    .A_N(_02408_));
 sg13g2_mux2_2 _07836_ (.A0(\cpu.PCreg0[5] ),
    .A1(\cpu.PCreg1[5] ),
    .S(net3636),
    .X(\cpu.PC[5] ));
 sg13g2_xnor2_1 _07837_ (.Y(_02415_),
    .A(_01664_),
    .B(_01871_));
 sg13g2_xor2_1 _07838_ (.B(_02415_),
    .A(_01978_),
    .X(_02416_));
 sg13g2_mux2_1 _07839_ (.A0(\cpu.PC[5] ),
    .A1(_02416_),
    .S(net3405),
    .X(_02417_));
 sg13g2_inv_1 _07840_ (.Y(_02418_),
    .A(net3128));
 sg13g2_nor2_1 _07841_ (.A(_02414_),
    .B(net3128),
    .Y(_02419_));
 sg13g2_xnor2_1 _07842_ (.Y(_02420_),
    .A(_01931_),
    .B(_01973_));
 sg13g2_mux2_2 _07843_ (.A0(\cpu.PCreg0[2] ),
    .A1(\cpu.PCreg1[2] ),
    .S(net3637),
    .X(\cpu.PC[2] ));
 sg13g2_mux2_1 _07844_ (.A0(_02420_),
    .A1(\cpu.PC[2] ),
    .S(net3406),
    .X(_02421_));
 sg13g2_nor3_1 _07845_ (.A(_02414_),
    .B(net3128),
    .C(net3142),
    .Y(_02422_));
 sg13g2_nand2_1 _07846_ (.Y(_02423_),
    .A(net3098),
    .B(_02422_));
 sg13g2_nor3_1 _07847_ (.A(\uart0.rxvalid ),
    .B(net3450),
    .C(_02423_),
    .Y(_02424_));
 sg13g2_nor4_2 _07848_ (.A(\uart0.txbitcnt[3] ),
    .B(\uart0.txbitcnt[2] ),
    .C(\uart0.txbitcnt[1] ),
    .Y(_02425_),
    .D(\uart0.txbitcnt[0] ));
 sg13g2_nor2_1 _07849_ (.A(\cpu.IR[6] ),
    .B(_01696_),
    .Y(_02426_));
 sg13g2_nand2b_1 _07850_ (.Y(_02427_),
    .B(\cpu.IR[4] ),
    .A_N(\cpu.IR[6] ));
 sg13g2_nand3_1 _07851_ (.B(\cpu.IR[1] ),
    .C(\cpu.IR[0] ),
    .A(\cpu.IR[2] ),
    .Y(_02428_));
 sg13g2_nor2_1 _07852_ (.A(_01759_),
    .B(_02428_),
    .Y(_02429_));
 sg13g2_nor3_1 _07853_ (.A(_01759_),
    .B(_02427_),
    .C(_02428_),
    .Y(_02430_));
 sg13g2_nand2_2 _07854_ (.Y(_02431_),
    .A(_02426_),
    .B(_02429_));
 sg13g2_and2_2 _07855_ (.A(_01947_),
    .B(net3394),
    .X(_02432_));
 sg13g2_nand2_1 _07856_ (.Y(_02433_),
    .A(_01947_),
    .B(net3394));
 sg13g2_nand2b_2 _07857_ (.Y(_02434_),
    .B(\cpu.IR[5] ),
    .A_N(_00547_));
 sg13g2_nor3_2 _07858_ (.A(\cpu.IR[4] ),
    .B(_01760_),
    .C(_02434_),
    .Y(_02435_));
 sg13g2_nor2_2 _07859_ (.A(_01760_),
    .B(_02427_),
    .Y(_02436_));
 sg13g2_nand2b_2 _07860_ (.Y(_02437_),
    .B(_02426_),
    .A_N(_01760_));
 sg13g2_nand2_1 _07861_ (.Y(_02438_),
    .A(net3696),
    .B(_00552_));
 sg13g2_nand2b_1 _07862_ (.Y(_02439_),
    .B(\cpu.IR[5] ),
    .A_N(_00562_));
 sg13g2_a21oi_1 _07863_ (.A1(_02438_),
    .A2(_02439_),
    .Y(_02440_),
    .B1(_02437_));
 sg13g2_nor2_1 _07864_ (.A(_02435_),
    .B(_02440_),
    .Y(_02441_));
 sg13g2_or2_1 _07865_ (.X(_02442_),
    .B(_02440_),
    .A(_02435_));
 sg13g2_a21oi_1 _07866_ (.A1(\cpu.IR[5] ),
    .A2(_02436_),
    .Y(_02443_),
    .B1(_02435_));
 sg13g2_a21o_2 _07867_ (.A2(_02436_),
    .A1(\cpu.IR[5] ),
    .B1(_02435_),
    .X(_02444_));
 sg13g2_and2_1 _07868_ (.A(\cpu.IR[21] ),
    .B(net3701),
    .X(_02445_));
 sg13g2_nand2_1 _07869_ (.Y(_02446_),
    .A(\cpu.IR[21] ),
    .B(net3700));
 sg13g2_and2_1 _07870_ (.A(net3646),
    .B(net3702),
    .X(_02447_));
 sg13g2_nand2_1 _07871_ (.Y(_02448_),
    .A(net3645),
    .B(net3700));
 sg13g2_and2_1 _07872_ (.A(\cpu.IR[22] ),
    .B(net3700),
    .X(_02449_));
 sg13g2_nand2_1 _07873_ (.Y(_02450_),
    .A(\cpu.IR[22] ),
    .B(net3700));
 sg13g2_mux4_1 _07874_ (.S0(net3480),
    .A0(_01680_),
    .A1(_01681_),
    .A2(_01682_),
    .A3(_01683_),
    .S1(net3532),
    .X(_02451_));
 sg13g2_and2_2 _07875_ (.A(\cpu.IR[23] ),
    .B(net3701),
    .X(_02452_));
 sg13g2_nand2_1 _07876_ (.Y(_02453_),
    .A(\cpu.IR[23] ),
    .B(net3700));
 sg13g2_a21oi_1 _07877_ (.A1(_01684_),
    .A2(net3480),
    .Y(_02454_),
    .B1(net3533));
 sg13g2_o21ai_1 _07878_ (.B1(_02454_),
    .Y(_02455_),
    .A1(_00540_),
    .A2(net3480));
 sg13g2_mux2_1 _07879_ (.A0(_00188_),
    .A1(_00316_),
    .S(net3480),
    .X(_02456_));
 sg13g2_a21oi_1 _07880_ (.A1(net3533),
    .A2(_02456_),
    .Y(_02457_),
    .B1(net3467));
 sg13g2_a221oi_1 _07881_ (.B2(_02457_),
    .C1(net3462),
    .B1(_02455_),
    .A1(net3467),
    .Y(_02458_),
    .A2(_02451_));
 sg13g2_nor2_2 _07882_ (.A(\cpu.IR[23] ),
    .B(net3467),
    .Y(_02459_));
 sg13g2_mux4_1 _07883_ (.S0(net3481),
    .A0(_00252_),
    .A1(_00122_),
    .A2(_00412_),
    .A3(_00284_),
    .S1(net3532),
    .X(_02460_));
 sg13g2_and2_1 _07884_ (.A(net3431),
    .B(_02460_),
    .X(_02461_));
 sg13g2_nor2_1 _07885_ (.A(net3471),
    .B(_02452_),
    .Y(_02462_));
 sg13g2_nand2_2 _07886_ (.Y(_02463_),
    .A(net3465),
    .B(net3461));
 sg13g2_o21ai_1 _07887_ (.B1(net3518),
    .Y(_02464_),
    .A1(_00508_),
    .A2(net3481));
 sg13g2_nor2_1 _07888_ (.A(_00090_),
    .B(net3481),
    .Y(_02465_));
 sg13g2_o21ai_1 _07889_ (.B1(net3532),
    .Y(_02466_),
    .A1(_00380_),
    .A2(net3646));
 sg13g2_o21ai_1 _07890_ (.B1(_02464_),
    .Y(_02467_),
    .A1(_02465_),
    .A2(_02466_));
 sg13g2_a21o_1 _07891_ (.A2(_02467_),
    .A1(net3429),
    .B1(_02461_),
    .X(_02468_));
 sg13g2_nor2_2 _07892_ (.A(_02458_),
    .B(_02468_),
    .Y(_02469_));
 sg13g2_or3_2 _07893_ (.A(net3370),
    .B(_02458_),
    .C(_02468_),
    .X(_02470_));
 sg13g2_nor4_1 _07894_ (.A(\cpu.IR[4] ),
    .B(_01759_),
    .C(_02428_),
    .D(_02434_),
    .Y(_02471_));
 sg13g2_nand3b_1 _07895_ (.B(_01696_),
    .C(_02429_),
    .Y(_02472_),
    .A_N(_02434_));
 sg13g2_or2_2 _07896_ (.X(_02473_),
    .B(net3423),
    .A(_01762_));
 sg13g2_a22oi_1 _07897_ (.Y(_02474_),
    .B1(_02473_),
    .B2(\cpu.IR[21] ),
    .A2(net3451),
    .A1(\cpu.Bimm[1] ));
 sg13g2_and2_1 _07898_ (.A(_02470_),
    .B(_02474_),
    .X(_02475_));
 sg13g2_nand3_1 _07899_ (.B(_02470_),
    .C(_02474_),
    .A(net3335),
    .Y(_02476_));
 sg13g2_a21o_1 _07900_ (.A2(_02474_),
    .A1(_02470_),
    .B1(net3335),
    .X(_02477_));
 sg13g2_nand2_1 _07901_ (.Y(_02478_),
    .A(_02476_),
    .B(_02477_));
 sg13g2_nand3_1 _07902_ (.B(_02476_),
    .C(_02477_),
    .A(_02432_),
    .Y(_02479_));
 sg13g2_a21oi_1 _07903_ (.A1(_02476_),
    .A2(_02477_),
    .Y(_02480_),
    .B1(_02432_));
 sg13g2_xnor2_1 _07904_ (.Y(_02481_),
    .A(_02432_),
    .B(_02478_));
 sg13g2_nor3_2 _07905_ (.A(net3538),
    .B(net3512),
    .C(_02463_),
    .Y(_02482_));
 sg13g2_nand3_1 _07906_ (.B(net3491),
    .C(net3428),
    .A(net3522),
    .Y(_02483_));
 sg13g2_nand2b_1 _07907_ (.Y(_02484_),
    .B(net3511),
    .A_N(\cpu.regs[13][0] ));
 sg13g2_nand2b_1 _07908_ (.Y(_02485_),
    .B(net3645),
    .A_N(\cpu.regs[15][0] ));
 sg13g2_a21oi_1 _07909_ (.A1(_01687_),
    .A2(net3481),
    .Y(_02486_),
    .B1(net3532));
 sg13g2_a21oi_1 _07910_ (.A1(_01688_),
    .A2(net3481),
    .Y(_02487_),
    .B1(net3519));
 sg13g2_a221oi_1 _07911_ (.B2(_02485_),
    .C1(net3467),
    .B1(_02487_),
    .A1(_02484_),
    .Y(_02488_),
    .A2(_02486_));
 sg13g2_mux4_1 _07912_ (.S0(net3511),
    .A0(\cpu.regs[8][0] ),
    .A1(\cpu.regs[9][0] ),
    .A2(\cpu.regs[10][0] ),
    .A3(\cpu.regs[11][0] ),
    .S1(net3532),
    .X(_02489_));
 sg13g2_o21ai_1 _07913_ (.B1(_02452_),
    .Y(_02490_),
    .A1(net3472),
    .A2(_02489_));
 sg13g2_or2_1 _07914_ (.X(_02491_),
    .B(_02490_),
    .A(_02488_));
 sg13g2_nor2_1 _07915_ (.A(\cpu.regs[3][0] ),
    .B(net3478),
    .Y(_02492_));
 sg13g2_mux4_1 _07916_ (.S0(net3516),
    .A0(\cpu.regs[4][0] ),
    .A1(\cpu.regs[5][0] ),
    .A2(\cpu.regs[6][0] ),
    .A3(\cpu.regs[7][0] ),
    .S1(net3531),
    .X(_02493_));
 sg13g2_nand2_1 _07917_ (.Y(_02494_),
    .A(\cpu.regs[1][0] ),
    .B(net3519));
 sg13g2_o21ai_1 _07918_ (.B1(net3531),
    .Y(_02495_),
    .A1(\cpu.regs[2][0] ),
    .A2(net3645));
 sg13g2_o21ai_1 _07919_ (.B1(_02494_),
    .Y(_02496_),
    .A1(_02492_),
    .A2(_02495_));
 sg13g2_a22oi_1 _07920_ (.Y(_02497_),
    .B1(_02496_),
    .B2(net3429),
    .A2(_02493_),
    .A1(net3430));
 sg13g2_a21oi_2 _07921_ (.B1(net3386),
    .Y(_02498_),
    .A2(_02497_),
    .A1(_02491_));
 sg13g2_and2_1 _07922_ (.A(\cpu.Bimm[11] ),
    .B(net3451),
    .X(_02499_));
 sg13g2_a221oi_1 _07923_ (.B2(net3368),
    .C1(_02499_),
    .B1(_02498_),
    .A1(net3645),
    .Y(_02500_),
    .A2(_02473_));
 sg13g2_and2_2 _07924_ (.A(_01968_),
    .B(net3393),
    .X(_02501_));
 sg13g2_nand2_2 _07925_ (.Y(_02502_),
    .A(_01968_),
    .B(net3393));
 sg13g2_mux2_1 _07926_ (.A0(_02502_),
    .A1(net3336),
    .S(net3289),
    .X(_02503_));
 sg13g2_xnor2_1 _07927_ (.Y(_02504_),
    .A(_02481_),
    .B(_02503_));
 sg13g2_inv_2 _07928_ (.Y(_02505_),
    .A(net3138));
 sg13g2_nor2_2 _07929_ (.A(net3695),
    .B(net3134),
    .Y(_02506_));
 sg13g2_nand2_1 _07930_ (.Y(_02507_),
    .A(net3625),
    .B(net3138));
 sg13g2_xnor2_1 _07931_ (.Y(_02508_),
    .A(net3289),
    .B(_02501_));
 sg13g2_nor2_2 _07932_ (.A(net3699),
    .B(net3698),
    .Y(_02509_));
 sg13g2_nand2_2 _07933_ (.Y(_02510_),
    .A(_01697_),
    .B(net3624));
 sg13g2_and2_1 _07934_ (.A(net3236),
    .B(net3459),
    .X(_02511_));
 sg13g2_nand2_2 _07935_ (.Y(_02512_),
    .A(net3236),
    .B(_02509_));
 sg13g2_nor2_2 _07936_ (.A(_01697_),
    .B(net3695),
    .Y(_02513_));
 sg13g2_nand2_2 _07937_ (.Y(_02514_),
    .A(net3699),
    .B(net3625));
 sg13g2_nor2_2 _07938_ (.A(net3134),
    .B(_02514_),
    .Y(_02515_));
 sg13g2_nor2_1 _07939_ (.A(net3135),
    .B(net3231),
    .Y(_02516_));
 sg13g2_nor2_2 _07940_ (.A(_02506_),
    .B(_02511_),
    .Y(_02517_));
 sg13g2_nand2_2 _07941_ (.Y(_02518_),
    .A(_02507_),
    .B(_02512_));
 sg13g2_and2_1 _07942_ (.A(net3450),
    .B(_02517_),
    .X(_02519_));
 sg13g2_nand2_1 _07943_ (.Y(_02520_),
    .A(net3450),
    .B(_02517_));
 sg13g2_nor2_1 _07944_ (.A(_02423_),
    .B(_02520_),
    .Y(_02521_));
 sg13g2_nor3_1 _07945_ (.A(_02423_),
    .B(_02425_),
    .C(_02520_),
    .Y(_02522_));
 sg13g2_nor3_1 _07946_ (.A(_01540_),
    .B(net3450),
    .C(_02423_),
    .Y(_02523_));
 sg13g2_nand3b_1 _07947_ (.B(net3739),
    .C(\uart0.rxoverr ),
    .Y(_02524_),
    .A_N(_02523_));
 sg13g2_o21ai_1 _07948_ (.B1(_02524_),
    .Y(_01531_),
    .A1(_01540_),
    .A2(net3739));
 sg13g2_o21ai_1 _07949_ (.B1(net3739),
    .Y(_01530_),
    .A1(_01540_),
    .A2(_02523_));
 sg13g2_mux2_1 _07950_ (.A0(\uart0.urxsh[9] ),
    .A1(\uart0.urxbuffer[8] ),
    .S(net3738),
    .X(_01529_));
 sg13g2_mux2_1 _07951_ (.A0(\uart0.urxsh[8] ),
    .A1(\uart0.q[7] ),
    .S(net3738),
    .X(_01528_));
 sg13g2_mux2_1 _07952_ (.A0(\uart0.urxsh[7] ),
    .A1(\uart0.q[6] ),
    .S(net3738),
    .X(_01527_));
 sg13g2_mux2_1 _07953_ (.A0(\uart0.urxsh[6] ),
    .A1(\uart0.q[5] ),
    .S(net3738),
    .X(_01526_));
 sg13g2_mux2_1 _07954_ (.A0(\uart0.urxsh[5] ),
    .A1(\uart0.q[4] ),
    .S(net3738),
    .X(_01525_));
 sg13g2_mux2_1 _07955_ (.A0(\uart0.urxsh[4] ),
    .A1(\uart0.q[3] ),
    .S(net3738),
    .X(_01524_));
 sg13g2_nor2_1 _07956_ (.A(net3739),
    .B(\uart0.urxsh[3] ),
    .Y(_02525_));
 sg13g2_a21oi_1 _07957_ (.A1(net3739),
    .A2(_01541_),
    .Y(_01523_),
    .B1(_02525_));
 sg13g2_mux2_1 _07958_ (.A0(\uart0.urxsh[2] ),
    .A1(\uart0.q[1] ),
    .S(net3739),
    .X(_01522_));
 sg13g2_mux2_1 _07959_ (.A0(\uart0.urxsh[1] ),
    .A1(\uart0.q[0] ),
    .S(net3739),
    .X(_01521_));
 sg13g2_nand3b_1 _07960_ (.B(_02425_),
    .C(_02521_),
    .Y(_02526_),
    .A_N(_02424_));
 sg13g2_nor3_1 _07961_ (.A(\uart0.txdiv[3] ),
    .B(\uart0.txdiv[2] ),
    .C(\uart0.txdiv[4] ),
    .Y(_02527_));
 sg13g2_nand4_1 _07962_ (.B(\uart0.txdiv[1] ),
    .C(\uart0.txdiv[5] ),
    .A(_01701_),
    .Y(_02528_),
    .D(_02527_));
 sg13g2_nor2_1 _07963_ (.A(_02425_),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_inv_1 _07964_ (.Y(_02530_),
    .A(_02529_));
 sg13g2_or4_1 _07965_ (.A(\uart0.txbitcnt[2] ),
    .B(\uart0.txbitcnt[1] ),
    .C(\uart0.txbitcnt[0] ),
    .D(_02530_),
    .X(_02531_));
 sg13g2_nand2_1 _07966_ (.Y(_02532_),
    .A(\uart0.txbitcnt[3] ),
    .B(_02531_));
 sg13g2_nand2_1 _07967_ (.Y(_01520_),
    .A(net3050),
    .B(_02532_));
 sg13g2_nor3_1 _07968_ (.A(\uart0.txbitcnt[1] ),
    .B(\uart0.txbitcnt[0] ),
    .C(_02528_),
    .Y(_02533_));
 sg13g2_o21ai_1 _07969_ (.B1(_02531_),
    .Y(_01519_),
    .A1(_01542_),
    .A2(_02533_));
 sg13g2_a21oi_1 _07970_ (.A1(net3050),
    .A2(_02530_),
    .Y(_02534_),
    .B1(\uart0.txbitcnt[0] ));
 sg13g2_xor2_1 _07971_ (.B(_02534_),
    .A(\uart0.txbitcnt[1] ),
    .X(_01518_));
 sg13g2_and3_1 _07972_ (.X(_02535_),
    .A(\uart0.txbitcnt[0] ),
    .B(net3050),
    .C(_02528_));
 sg13g2_a21o_1 _07973_ (.A2(_02534_),
    .A1(net3050),
    .B1(_02535_),
    .X(_01517_));
 sg13g2_nor2_1 _07974_ (.A(\uart0.rxdiv[0] ),
    .B(\uart0.rxdiv[1] ),
    .Y(_02536_));
 sg13g2_nor3_1 _07975_ (.A(\uart0.rxdiv[3] ),
    .B(\uart0.rxdiv[2] ),
    .C(\uart0.rxdiv[5] ),
    .Y(_02537_));
 sg13g2_nand3_1 _07976_ (.B(_02536_),
    .C(_02537_),
    .A(\uart0.rxdiv[4] ),
    .Y(_02538_));
 sg13g2_and2_1 _07977_ (.A(net3738),
    .B(_02538_),
    .X(_02539_));
 sg13g2_nand2_1 _07978_ (.Y(_02540_),
    .A(_00590_),
    .B(net3417));
 sg13g2_nand4_1 _07979_ (.B(\uart0.rxdiv[4] ),
    .C(_02536_),
    .A(net3738),
    .Y(_02541_),
    .D(_02537_));
 sg13g2_o21ai_1 _07980_ (.B1(_02540_),
    .Y(_01516_),
    .A1(\uart0.rxreg[1] ),
    .A2(net3458));
 sg13g2_nand2_1 _07981_ (.Y(_02542_),
    .A(_00589_),
    .B(net3417));
 sg13g2_o21ai_1 _07982_ (.B1(_02542_),
    .Y(_01515_),
    .A1(\uart0.urxsh[9] ),
    .A2(net3458));
 sg13g2_nand2_1 _07983_ (.Y(_02543_),
    .A(_00588_),
    .B(net3417));
 sg13g2_o21ai_1 _07984_ (.B1(_02543_),
    .Y(_01514_),
    .A1(\uart0.urxsh[8] ),
    .A2(net3458));
 sg13g2_nand2_1 _07985_ (.Y(_02544_),
    .A(_00587_),
    .B(net3417));
 sg13g2_o21ai_1 _07986_ (.B1(_02544_),
    .Y(_01513_),
    .A1(\uart0.urxsh[7] ),
    .A2(net3458));
 sg13g2_nand2_1 _07987_ (.Y(_02545_),
    .A(_00586_),
    .B(net3417));
 sg13g2_o21ai_1 _07988_ (.B1(_02545_),
    .Y(_01512_),
    .A1(\uart0.urxsh[6] ),
    .A2(net3458));
 sg13g2_nand2_1 _07989_ (.Y(_02546_),
    .A(_00585_),
    .B(net3417));
 sg13g2_o21ai_1 _07990_ (.B1(_02546_),
    .Y(_01511_),
    .A1(\uart0.urxsh[5] ),
    .A2(net3458));
 sg13g2_nand2_1 _07991_ (.Y(_02547_),
    .A(_00584_),
    .B(net3417));
 sg13g2_o21ai_1 _07992_ (.B1(_02547_),
    .Y(_01510_),
    .A1(\uart0.urxsh[4] ),
    .A2(net3458));
 sg13g2_nand2_1 _07993_ (.Y(_02548_),
    .A(_00583_),
    .B(_02539_));
 sg13g2_o21ai_1 _07994_ (.B1(_02548_),
    .Y(_01509_),
    .A1(\uart0.urxsh[3] ),
    .A2(_02541_));
 sg13g2_nand2_1 _07995_ (.Y(_02549_),
    .A(_00582_),
    .B(net3417));
 sg13g2_o21ai_1 _07996_ (.B1(_02549_),
    .Y(_01508_),
    .A1(\uart0.urxsh[2] ),
    .A2(net3458));
 sg13g2_nor2_1 _07997_ (.A(\uart0.urxsh[1] ),
    .B(_02541_),
    .Y(_00691_));
 sg13g2_nand2_1 _07998_ (.Y(_02550_),
    .A(_01700_),
    .B(net3926));
 sg13g2_nand3_1 _07999_ (.B(\jtag0.tapst[1] ),
    .C(net3926),
    .A(net3927),
    .Y(_02551_));
 sg13g2_nor2_1 _08000_ (.A(\jtag0.tapst[3] ),
    .B(_02551_),
    .Y(_02552_));
 sg13g2_nor2_1 _08001_ (.A(\bsq[29] ),
    .B(net3906),
    .Y(_02553_));
 sg13g2_a21oi_1 _08002_ (.A1(_01543_),
    .A2(net3906),
    .Y(_01345_),
    .B1(_02553_));
 sg13g2_nor2_1 _08003_ (.A(\bsq[28] ),
    .B(net3906),
    .Y(_02554_));
 sg13g2_a21oi_1 _08004_ (.A1(_01544_),
    .A2(net3906),
    .Y(_01344_),
    .B1(_02554_));
 sg13g2_nor2_1 _08005_ (.A(\bsq[27] ),
    .B(net3906),
    .Y(_02555_));
 sg13g2_a21oi_1 _08006_ (.A1(_01545_),
    .A2(net3906),
    .Y(_01343_),
    .B1(_02555_));
 sg13g2_mux2_1 _08007_ (.A0(\bsq[26] ),
    .A1(\jtag0.bssh[26] ),
    .S(net3906),
    .X(_01342_));
 sg13g2_mux2_1 _08008_ (.A0(\bsq[25] ),
    .A1(\jtag0.bssh[25] ),
    .S(net3908),
    .X(_01341_));
 sg13g2_nor2_1 _08009_ (.A(\bsq[24] ),
    .B(net3909),
    .Y(_02556_));
 sg13g2_a21oi_1 _08010_ (.A1(_01546_),
    .A2(net3909),
    .Y(_01340_),
    .B1(_02556_));
 sg13g2_nor2_1 _08011_ (.A(\bsq[23] ),
    .B(net3908),
    .Y(_02557_));
 sg13g2_a21oi_1 _08012_ (.A1(_01547_),
    .A2(net3908),
    .Y(_01339_),
    .B1(_02557_));
 sg13g2_nor2_1 _08013_ (.A(\bsq[22] ),
    .B(net3905),
    .Y(_02558_));
 sg13g2_a21oi_1 _08014_ (.A1(_01548_),
    .A2(net3904),
    .Y(_01338_),
    .B1(_02558_));
 sg13g2_nor2_1 _08015_ (.A(\bsq[21] ),
    .B(net3905),
    .Y(_02559_));
 sg13g2_a21oi_1 _08016_ (.A1(_01549_),
    .A2(net3904),
    .Y(_01337_),
    .B1(_02559_));
 sg13g2_mux2_1 _08017_ (.A0(\bsq[20] ),
    .A1(\jtag0.bssh[20] ),
    .S(net3906),
    .X(_01336_));
 sg13g2_mux2_1 _08018_ (.A0(\bsq[19] ),
    .A1(\jtag0.bssh[19] ),
    .S(net3907),
    .X(_01335_));
 sg13g2_nor2_1 _08019_ (.A(\bsq[18] ),
    .B(net3907),
    .Y(_02560_));
 sg13g2_a21oi_1 _08020_ (.A1(_01550_),
    .A2(net3907),
    .Y(_01334_),
    .B1(_02560_));
 sg13g2_nor2_1 _08021_ (.A(\bsq[17] ),
    .B(net3905),
    .Y(_02561_));
 sg13g2_a21oi_1 _08022_ (.A1(_01551_),
    .A2(net3905),
    .Y(_01333_),
    .B1(_02561_));
 sg13g2_nor2_1 _08023_ (.A(\bsq[16] ),
    .B(net3908),
    .Y(_02562_));
 sg13g2_a21oi_1 _08024_ (.A1(_01552_),
    .A2(net3908),
    .Y(_01332_),
    .B1(_02562_));
 sg13g2_nor2_1 _08025_ (.A(\bsq[15] ),
    .B(net3908),
    .Y(_02563_));
 sg13g2_a21oi_1 _08026_ (.A1(_01553_),
    .A2(net3908),
    .Y(_01331_),
    .B1(_02563_));
 sg13g2_mux2_1 _08027_ (.A0(\bsq[14] ),
    .A1(\jtag0.bssh[14] ),
    .S(net3910),
    .X(_01330_));
 sg13g2_mux2_1 _08028_ (.A0(\bsq[13] ),
    .A1(\jtag0.bssh[13] ),
    .S(net3910),
    .X(_01329_));
 sg13g2_mux2_1 _08029_ (.A0(\bsq[12] ),
    .A1(\jtag0.bssh[12] ),
    .S(net3908),
    .X(_01328_));
 sg13g2_mux2_1 _08030_ (.A0(\bsq[11] ),
    .A1(\jtag0.bssh[11] ),
    .S(net3909),
    .X(_01327_));
 sg13g2_mux2_1 _08031_ (.A0(\bsq[10] ),
    .A1(\jtag0.bssh[10] ),
    .S(net3909),
    .X(_01326_));
 sg13g2_mux2_1 _08032_ (.A0(\bsq[9] ),
    .A1(\jtag0.bssh[9] ),
    .S(net3910),
    .X(_01325_));
 sg13g2_mux2_1 _08033_ (.A0(\bsq[8] ),
    .A1(\jtag0.bssh[8] ),
    .S(net3909),
    .X(_01324_));
 sg13g2_mux2_1 _08034_ (.A0(\bsq[7] ),
    .A1(\jtag0.bssh[7] ),
    .S(net3909),
    .X(_01323_));
 sg13g2_mux2_1 _08035_ (.A0(\bsq[6] ),
    .A1(\jtag0.bssh[6] ),
    .S(net3909),
    .X(_01322_));
 sg13g2_mux2_1 _08036_ (.A0(\bsq[5] ),
    .A1(\jtag0.bssh[5] ),
    .S(net3909),
    .X(_01321_));
 sg13g2_mux2_1 _08037_ (.A0(\bsq[4] ),
    .A1(\jtag0.bssh[4] ),
    .S(net3904),
    .X(_01320_));
 sg13g2_mux2_1 _08038_ (.A0(\bsq[3] ),
    .A1(\jtag0.bssh[3] ),
    .S(net3904),
    .X(_01319_));
 sg13g2_mux2_1 _08039_ (.A0(\bsq[2] ),
    .A1(\jtag0.bssh[2] ),
    .S(net3904),
    .X(_01318_));
 sg13g2_mux2_1 _08040_ (.A0(\bsq[1] ),
    .A1(\jtag0.bssh[1] ),
    .S(net3904),
    .X(_01317_));
 sg13g2_nor2_1 _08041_ (.A(\bsq[0] ),
    .B(net3904),
    .Y(_02564_));
 sg13g2_a21oi_1 _08042_ (.A1(_01554_),
    .A2(net3904),
    .Y(_01316_),
    .B1(_02564_));
 sg13g2_nand2_1 _08043_ (.Y(_02565_),
    .A(\jtag0.ir[1] ),
    .B(_00125_));
 sg13g2_inv_1 _08044_ (.Y(_00003_),
    .A(_02565_));
 sg13g2_nor2_1 _08045_ (.A(_01573_),
    .B(_02565_),
    .Y(_02566_));
 sg13g2_nand2_1 _08046_ (.Y(_02567_),
    .A(\jtag0.ir[0] ),
    .B(_00003_));
 sg13g2_nand4_1 _08047_ (.B(_02397_),
    .C(_02398_),
    .A(_02396_),
    .Y(_02568_),
    .D(_02400_));
 sg13g2_nor3_1 _08048_ (.A(_01767_),
    .B(_02387_),
    .C(_02568_),
    .Y(_02569_));
 sg13g2_inv_2 _08049_ (.Y(_02570_),
    .A(net3096));
 sg13g2_nand2_1 _08050_ (.Y(_02571_),
    .A(net3925),
    .B(net3450));
 sg13g2_nor2_1 _08051_ (.A(\ckd[1] ),
    .B(_02519_),
    .Y(_02572_));
 sg13g2_o21ai_1 _08052_ (.B1(_02572_),
    .Y(_02573_),
    .A1(_02515_),
    .A2(_02571_));
 sg13g2_nor2_2 _08053_ (.A(_01707_),
    .B(\ckd[1] ),
    .Y(_02574_));
 sg13g2_nor2b_1 _08054_ (.A(net3925),
    .B_N(\ckd[1] ),
    .Y(_02575_));
 sg13g2_o21ai_1 _08055_ (.B1(net3235),
    .Y(_02576_),
    .A1(\ckd[1] ),
    .A2(net3134));
 sg13g2_a22oi_1 _08056_ (.Y(_02577_),
    .B1(_02576_),
    .B2(net3925),
    .A2(_02575_),
    .A1(net3235));
 sg13g2_nor2_1 _08057_ (.A(_02510_),
    .B(_02577_),
    .Y(_02578_));
 sg13g2_nand2_1 _08058_ (.Y(_02579_),
    .A(net3698),
    .B(net3450));
 sg13g2_nand2_1 _08059_ (.Y(_02580_),
    .A(\ckd[1] ),
    .B(_02579_));
 sg13g2_a21oi_1 _08060_ (.A1(net3450),
    .A2(net3139),
    .Y(_02581_),
    .B1(_02580_));
 sg13g2_mux2_1 _08061_ (.A0(clknet_1_1__leaf_clk),
    .A1(bsq1r),
    .S(net3929),
    .X(jclk));
 sg13g2_nor4_1 _08062_ (.A(net3923),
    .B(_02578_),
    .C(_02581_),
    .D(clknet_1_1__leaf_jclk),
    .Y(_02582_));
 sg13g2_nand3_1 _08063_ (.B(_02573_),
    .C(_02582_),
    .A(net3096),
    .Y(_02583_));
 sg13g2_mux2_1 _08064_ (.A0(clknet_1_1__leaf__02583_),
    .A1(\bsq[29] ),
    .S(net3930),
    .X(uo_out[7]));
 sg13g2_nor2_1 _08065_ (.A(net3900),
    .B(uo_out[7]),
    .Y(_02584_));
 sg13g2_nor2_2 _08066_ (.A(\jtag0.tapst[3] ),
    .B(net3926),
    .Y(_02585_));
 sg13g2_and2_2 _08067_ (.A(\jtag0.tapst[1] ),
    .B(_02585_),
    .X(_02586_));
 sg13g2_nand2_1 _08068_ (.Y(_02587_),
    .A(\jtag0.tapst[1] ),
    .B(_02585_));
 sg13g2_nor2_1 _08069_ (.A(net3928),
    .B(net3892),
    .Y(_02588_));
 sg13g2_nand2b_2 _08070_ (.Y(_02589_),
    .B(_02586_),
    .A_N(net3927));
 sg13g2_o21ai_1 _08071_ (.B1(net3729),
    .Y(_02590_),
    .A1(net3735),
    .A2(clknet_1_0__leaf__02583_));
 sg13g2_nor2b_1 _08072_ (.A(_01752_),
    .B_N(_02585_),
    .Y(_02591_));
 sg13g2_a22oi_1 _08073_ (.Y(_02592_),
    .B1(net3885),
    .B2(\jtag0.stdi ),
    .A2(net3892),
    .A1(\jtag0.bssh[29] ));
 sg13g2_o21ai_1 _08074_ (.B1(_02592_),
    .Y(_01315_),
    .A1(_02584_),
    .A2(_02590_));
 sg13g2_nor3_2 _08075_ (.A(net3919),
    .B(net3451),
    .C(_02570_),
    .Y(_02593_));
 sg13g2_nand2_1 _08076_ (.Y(_02594_),
    .A(\bsq[28] ),
    .B(net3930));
 sg13g2_o21ai_1 _08077_ (.B1(_02594_),
    .Y(net3049),
    .A1(net3930),
    .A2(_02593_));
 sg13g2_o21ai_1 _08078_ (.B1(net3730),
    .Y(_02595_),
    .A1(net3735),
    .A2(_02593_));
 sg13g2_a21oi_1 _08079_ (.A1(net3735),
    .A2(net3049),
    .Y(_02596_),
    .B1(_02595_));
 sg13g2_a221oi_1 _08080_ (.B2(_01543_),
    .C1(_02596_),
    .B1(net3885),
    .A1(_01544_),
    .Y(_01314_),
    .A2(net3892));
 sg13g2_nand2_2 _08081_ (.Y(_02597_),
    .A(\ckd[1] ),
    .B(net3096));
 sg13g2_nand2_1 _08082_ (.Y(_02598_),
    .A(\bsq[27] ),
    .B(net3931));
 sg13g2_o21ai_1 _08083_ (.B1(_02598_),
    .Y(uo_out[5]),
    .A1(net3933),
    .A2(_02597_));
 sg13g2_a21oi_1 _08084_ (.A1(net3901),
    .A2(_02597_),
    .Y(_02599_),
    .B1(_02589_));
 sg13g2_o21ai_1 _08085_ (.B1(_02599_),
    .Y(_02600_),
    .A1(net3900),
    .A2(uo_out[5]));
 sg13g2_a21oi_1 _08086_ (.A1(\jtag0.bssh[28] ),
    .A2(net3928),
    .Y(_02601_),
    .B1(net3892));
 sg13g2_a22oi_1 _08087_ (.Y(_01313_),
    .B1(_02600_),
    .B2(_02601_),
    .A2(net3892),
    .A1(_01545_));
 sg13g2_mux2_2 _08088_ (.A0(txd),
    .A1(\bsq[26] ),
    .S(net3930),
    .X(uo_out[4]));
 sg13g2_nor2_1 _08089_ (.A(txd),
    .B(net3735),
    .Y(_02602_));
 sg13g2_o21ai_1 _08090_ (.B1(net3730),
    .Y(_02603_),
    .A1(net3900),
    .A2(uo_out[4]));
 sg13g2_a22oi_1 _08091_ (.Y(_02604_),
    .B1(net3885),
    .B2(\jtag0.bssh[27] ),
    .A2(net3893),
    .A1(\jtag0.bssh[26] ));
 sg13g2_o21ai_1 _08092_ (.B1(_02604_),
    .Y(_01312_),
    .A1(_02602_),
    .A2(_02603_));
 sg13g2_nand2_1 _08093_ (.Y(_02605_),
    .A(\jtag0.bssh[25] ),
    .B(net3894));
 sg13g2_a21oi_1 _08094_ (.A1(\jtag0.bssh[26] ),
    .A2(_02586_),
    .Y(_02606_),
    .B1(net3730));
 sg13g2_nand2_1 _08095_ (.Y(_02607_),
    .A(\bsq[25] ),
    .B(net3932));
 sg13g2_nor3_1 _08096_ (.A(_01707_),
    .B(net3932),
    .C(_02570_),
    .Y(_02608_));
 sg13g2_inv_1 _08097_ (.Y(_02609_),
    .A(_02608_));
 sg13g2_o21ai_1 _08098_ (.B1(_02607_),
    .Y(uo_out[2]),
    .A1(\ckd[2] ),
    .A2(_02609_));
 sg13g2_nand3_1 _08099_ (.B(net3902),
    .C(net3096),
    .A(net3925),
    .Y(_02610_));
 sg13g2_o21ai_1 _08100_ (.B1(net3731),
    .Y(_02611_),
    .A1(\ckd[2] ),
    .A2(_02610_));
 sg13g2_a21oi_1 _08101_ (.A1(net3736),
    .A2(uo_out[2]),
    .Y(_02612_),
    .B1(_02611_));
 sg13g2_o21ai_1 _08102_ (.B1(_02605_),
    .Y(_01311_),
    .A1(_02606_),
    .A2(_02612_));
 sg13g2_nor3_2 _08103_ (.A(net3925),
    .B(\ckd[2] ),
    .C(_02570_),
    .Y(_02613_));
 sg13g2_mux2_1 _08104_ (.A0(_02613_),
    .A1(\bsq[24] ),
    .S(net3933),
    .X(uo_out[1]));
 sg13g2_o21ai_1 _08105_ (.B1(net3731),
    .Y(_02614_),
    .A1(net3901),
    .A2(uo_out[1]));
 sg13g2_inv_1 _08106_ (.Y(_02615_),
    .A(_02614_));
 sg13g2_o21ai_1 _08107_ (.B1(_02615_),
    .Y(_02616_),
    .A1(net3737),
    .A2(_02613_));
 sg13g2_a21oi_1 _08108_ (.A1(\jtag0.bssh[25] ),
    .A2(net3928),
    .Y(_02617_),
    .B1(net3894));
 sg13g2_a22oi_1 _08109_ (.Y(_01310_),
    .B1(_02616_),
    .B2(_02617_),
    .A2(net3895),
    .A1(_01546_));
 sg13g2_a21oi_1 _08110_ (.A1(\bsq[23] ),
    .A2(net3932),
    .Y(_02618_),
    .B1(_02608_));
 sg13g2_inv_1 _08111_ (.Y(uo_out[0]),
    .A(_02618_));
 sg13g2_o21ai_1 _08112_ (.B1(_02610_),
    .Y(_02619_),
    .A1(net3902),
    .A2(_02618_));
 sg13g2_nand2_1 _08113_ (.Y(_02620_),
    .A(\jtag0.bssh[24] ),
    .B(net3882));
 sg13g2_a22oi_1 _08114_ (.Y(_02621_),
    .B1(net3731),
    .B2(_02619_),
    .A2(net3897),
    .A1(\jtag0.bssh[23] ));
 sg13g2_nand2_1 _08115_ (.Y(_01309_),
    .A(_02620_),
    .B(_02621_));
 sg13g2_and2_2 _08116_ (.A(net3921),
    .B(_02574_),
    .X(_02622_));
 sg13g2_nand2_1 _08117_ (.Y(_02623_),
    .A(net3921),
    .B(_02574_));
 sg13g2_mux2_2 _08118_ (.A0(\cpu.PCreg0[17] ),
    .A1(\cpu.PCreg1[17] ),
    .S(net3629),
    .X(\cpu.PC[17] ));
 sg13g2_o21ai_1 _08119_ (.B1(_02622_),
    .Y(_02624_),
    .A1(net3401),
    .A2(\cpu.PC[17] ));
 sg13g2_a21oi_1 _08120_ (.A1(net3642),
    .A2(_02118_),
    .Y(_02625_),
    .B1(_02120_));
 sg13g2_nor2_1 _08121_ (.A(_02223_),
    .B(_02224_),
    .Y(_02626_));
 sg13g2_xnor2_1 _08122_ (.Y(_02627_),
    .A(_02625_),
    .B(_02626_));
 sg13g2_a21oi_1 _08123_ (.A1(net3401),
    .A2(_02627_),
    .Y(_02628_),
    .B1(_02624_));
 sg13g2_nand2_1 _08124_ (.Y(_02629_),
    .A(net3925),
    .B(\ckd[1] ));
 sg13g2_nor2_1 _08125_ (.A(net3923),
    .B(_02629_),
    .Y(_02630_));
 sg13g2_nor2_1 _08126_ (.A(_00126_),
    .B(net3474),
    .Y(_02631_));
 sg13g2_o21ai_1 _08127_ (.B1(net3520),
    .Y(_02632_),
    .A1(_00190_),
    .A2(net3511));
 sg13g2_mux2_1 _08128_ (.A0(_00446_),
    .A1(_00318_),
    .S(net3475),
    .X(_02633_));
 sg13g2_o21ai_1 _08129_ (.B1(net3465),
    .Y(_02634_),
    .A1(_02631_),
    .A2(_02632_));
 sg13g2_a21oi_1 _08130_ (.A1(net3529),
    .A2(_02633_),
    .Y(_02635_),
    .B1(_02634_));
 sg13g2_nor2_1 _08131_ (.A(_00510_),
    .B(net3485),
    .Y(_02636_));
 sg13g2_o21ai_1 _08132_ (.B1(net3521),
    .Y(_02637_),
    .A1(_00414_),
    .A2(net3512));
 sg13g2_mux2_1 _08133_ (.A0(_00158_),
    .A1(_00286_),
    .S(net3485),
    .X(_02638_));
 sg13g2_o21ai_1 _08134_ (.B1(net3469),
    .Y(_02639_),
    .A1(_02636_),
    .A2(_02637_));
 sg13g2_a21oi_2 _08135_ (.B1(_02639_),
    .Y(_02640_),
    .A2(_02638_),
    .A1(net3537));
 sg13g2_nor3_1 _08136_ (.A(net3461),
    .B(_02635_),
    .C(_02640_),
    .Y(_02641_));
 sg13g2_mux4_1 _08137_ (.S0(net3477),
    .A0(_00222_),
    .A1(_00092_),
    .A2(_00382_),
    .A3(_00254_),
    .S1(net3530),
    .X(_02642_));
 sg13g2_nor2_1 _08138_ (.A(_00060_),
    .B(net3475),
    .Y(_02643_));
 sg13g2_o21ai_1 _08139_ (.B1(net3529),
    .Y(_02644_),
    .A1(net3647),
    .A2(_00350_));
 sg13g2_o21ai_1 _08140_ (.B1(net3517),
    .Y(_02645_),
    .A1(_00478_),
    .A2(net3475));
 sg13g2_o21ai_1 _08141_ (.B1(_02645_),
    .Y(_02646_),
    .A1(_02643_),
    .A2(_02644_));
 sg13g2_a221oi_1 _08142_ (.B2(net3426),
    .C1(_02641_),
    .B1(_02646_),
    .A1(net3430),
    .Y(_02647_),
    .A2(_02642_));
 sg13g2_nand2b_1 _08143_ (.Y(_02648_),
    .B(net3515),
    .A_N(_00150_));
 sg13g2_a21oi_1 _08144_ (.A1(_01645_),
    .A2(net3507),
    .Y(_02649_),
    .B1(net3551));
 sg13g2_mux2_1 _08145_ (.A0(_00470_),
    .A1(_00342_),
    .S(net3501),
    .X(_02650_));
 sg13g2_a221oi_1 _08146_ (.B2(net3551),
    .C1(net3473),
    .B1(_02650_),
    .A1(_02648_),
    .Y(_02651_),
    .A2(_02649_));
 sg13g2_mux2_1 _08147_ (.A0(_00534_),
    .A1(_00438_),
    .S(net3507),
    .X(_02652_));
 sg13g2_nand2_1 _08148_ (.Y(_02653_),
    .A(_01649_),
    .B(net3650));
 sg13g2_a21oi_1 _08149_ (.A1(_01650_),
    .A2(net3507),
    .Y(_02654_),
    .B1(net3526));
 sg13g2_a221oi_1 _08150_ (.B2(_02654_),
    .C1(net3466),
    .B1(_02653_),
    .A1(net3526),
    .Y(_02655_),
    .A2(_02652_));
 sg13g2_or3_1 _08151_ (.A(net3462),
    .B(_02651_),
    .C(_02655_),
    .X(_02656_));
 sg13g2_mux4_1 _08152_ (.S0(net3503),
    .A0(_00246_),
    .A1(_00116_),
    .A2(_00406_),
    .A3(_00278_),
    .S1(net3547),
    .X(_02657_));
 sg13g2_nor2_1 _08153_ (.A(_00084_),
    .B(net3503),
    .Y(_02658_));
 sg13g2_o21ai_1 _08154_ (.B1(net3547),
    .Y(_02659_),
    .A1(_00374_),
    .A2(net3651));
 sg13g2_o21ai_1 _08155_ (.B1(net3525),
    .Y(_02660_),
    .A1(_00502_),
    .A2(net3503));
 sg13g2_o21ai_1 _08156_ (.B1(_02660_),
    .Y(_02661_),
    .A1(_02658_),
    .A2(_02659_));
 sg13g2_a22oi_1 _08157_ (.Y(_02662_),
    .B1(_02661_),
    .B2(net3427),
    .A2(_02657_),
    .A1(net3433));
 sg13g2_and2_2 _08158_ (.A(_02656_),
    .B(_02662_),
    .X(_02663_));
 sg13g2_nand2b_1 _08159_ (.Y(_02664_),
    .B(net3515),
    .A_N(_00142_));
 sg13g2_a21oi_1 _08160_ (.A1(_01599_),
    .A2(net3499),
    .Y(_02665_),
    .B1(net3546));
 sg13g2_mux2_1 _08161_ (.A0(_00462_),
    .A1(_00334_),
    .S(net3499),
    .X(_02666_));
 sg13g2_a221oi_1 _08162_ (.B2(net3546),
    .C1(net3471),
    .B1(_02666_),
    .A1(_02664_),
    .Y(_02667_),
    .A2(_02665_));
 sg13g2_mux2_1 _08163_ (.A0(_00526_),
    .A1(_00430_),
    .S(net3499),
    .X(_02668_));
 sg13g2_nand2_1 _08164_ (.Y(_02669_),
    .A(_01603_),
    .B(net3650));
 sg13g2_a21oi_1 _08165_ (.A1(_01604_),
    .A2(net3499),
    .Y(_02670_),
    .B1(net3524));
 sg13g2_a221oi_1 _08166_ (.B2(_02670_),
    .C1(net3466),
    .B1(_02669_),
    .A1(net3524),
    .Y(_02671_),
    .A2(_02668_));
 sg13g2_or3_1 _08167_ (.A(net3463),
    .B(_02667_),
    .C(_02671_),
    .X(_02672_));
 sg13g2_mux4_1 _08168_ (.S0(net3500),
    .A0(_00238_),
    .A1(_00108_),
    .A2(_00398_),
    .A3(_00270_),
    .S1(net3546),
    .X(_02673_));
 sg13g2_nand2_1 _08169_ (.Y(_02674_),
    .A(net3433),
    .B(_02673_));
 sg13g2_nor2_1 _08170_ (.A(_00076_),
    .B(net3500),
    .Y(_02675_));
 sg13g2_o21ai_1 _08171_ (.B1(net3546),
    .Y(_02676_),
    .A1(_00366_),
    .A2(net3649));
 sg13g2_nand2_1 _08172_ (.Y(_02677_),
    .A(_00494_),
    .B(net3524));
 sg13g2_o21ai_1 _08173_ (.B1(_02677_),
    .Y(_02678_),
    .A1(_02675_),
    .A2(_02676_));
 sg13g2_nand2_1 _08174_ (.Y(_02679_),
    .A(net3427),
    .B(_02678_));
 sg13g2_nand4_1 _08175_ (.B(_02672_),
    .C(_02674_),
    .A(_02483_),
    .Y(_02680_),
    .D(_02679_));
 sg13g2_nor2_1 _08176_ (.A(net3232),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_a21oi_2 _08177_ (.B1(_02681_),
    .Y(_02682_),
    .A2(net3330),
    .A1(net3231));
 sg13g2_nor2_1 _08178_ (.A(net3130),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_a21oi_2 _08179_ (.B1(_02683_),
    .Y(_02684_),
    .A2(_02647_),
    .A1(net3130));
 sg13g2_inv_1 _08180_ (.Y(_02685_),
    .A(_02684_));
 sg13g2_nand2_1 _08181_ (.Y(_02686_),
    .A(\ckd[2] ),
    .B(_02575_));
 sg13g2_a21oi_1 _08182_ (.A1(_01722_),
    .A2(net3491),
    .Y(_02687_),
    .B1(net3540));
 sg13g2_o21ai_1 _08183_ (.B1(_02687_),
    .Y(_02688_),
    .A1(_00134_),
    .A2(net3491));
 sg13g2_mux2_1 _08184_ (.A0(_00454_),
    .A1(_00326_),
    .S(net3490),
    .X(_02689_));
 sg13g2_a21oi_1 _08185_ (.A1(net3545),
    .A2(_02689_),
    .Y(_02690_),
    .B1(net3469));
 sg13g2_a21oi_1 _08186_ (.A1(_01723_),
    .A2(net3491),
    .Y(_02691_),
    .B1(net3540));
 sg13g2_o21ai_1 _08187_ (.B1(_02691_),
    .Y(_02692_),
    .A1(_00518_),
    .A2(net3490));
 sg13g2_mux2_1 _08188_ (.A0(_00166_),
    .A1(_00294_),
    .S(net3491),
    .X(_02693_));
 sg13g2_a21oi_1 _08189_ (.A1(net3540),
    .A2(_02693_),
    .Y(_02694_),
    .B1(net3464));
 sg13g2_a221oi_1 _08190_ (.B2(_02694_),
    .C1(net3460),
    .B1(_02692_),
    .A1(_02688_),
    .Y(_02695_),
    .A2(_02690_));
 sg13g2_mux4_1 _08191_ (.S0(net3498),
    .A0(_00230_),
    .A1(_00100_),
    .A2(_00390_),
    .A3(_00262_),
    .S1(net3545),
    .X(_02696_));
 sg13g2_nor2_1 _08192_ (.A(_00068_),
    .B(net3492),
    .Y(_02697_));
 sg13g2_o21ai_1 _08193_ (.B1(net3540),
    .Y(_02698_),
    .A1(net3652),
    .A2(_00358_));
 sg13g2_o21ai_1 _08194_ (.B1(net3522),
    .Y(_02699_),
    .A1(_00486_),
    .A2(net3492));
 sg13g2_o21ai_1 _08195_ (.B1(_02699_),
    .Y(_02700_),
    .A1(_02697_),
    .A2(_02698_));
 sg13g2_a221oi_1 _08196_ (.B2(net3428),
    .C1(_02695_),
    .B1(_02700_),
    .A1(net3432),
    .Y(_02701_),
    .A2(_02696_));
 sg13g2_nor2b_2 _08197_ (.A(net3140),
    .B_N(_02701_),
    .Y(_02702_));
 sg13g2_a21oi_2 _08198_ (.B1(_02702_),
    .Y(_02703_),
    .A2(net3330),
    .A1(net3136));
 sg13g2_nor2_1 _08199_ (.A(net3725),
    .B(_02703_),
    .Y(_02704_));
 sg13g2_nand2_2 _08200_ (.Y(_02705_),
    .A(\ckd[2] ),
    .B(_02574_));
 sg13g2_nor2_1 _08201_ (.A(net3925),
    .B(\ckd[1] ),
    .Y(_02706_));
 sg13g2_and2_2 _08202_ (.A(\ckd[2] ),
    .B(_02706_),
    .X(_02707_));
 sg13g2_a221oi_1 _08203_ (.B2(net3330),
    .C1(_02704_),
    .B1(net3723),
    .A1(net3728),
    .Y(_02708_),
    .A2(_02685_));
 sg13g2_o21ai_1 _08204_ (.B1(_02708_),
    .Y(_02709_),
    .A1(_02682_),
    .A2(net3456));
 sg13g2_xnor2_1 _08205_ (.Y(_02710_),
    .A(_02018_),
    .B(_02034_));
 sg13g2_mux2_2 _08206_ (.A0(\cpu.PCreg0[9] ),
    .A1(\cpu.PCreg1[9] ),
    .S(net3635),
    .X(\cpu.PC[9] ));
 sg13g2_nand2_1 _08207_ (.Y(_02711_),
    .A(net927),
    .B(_02629_));
 sg13g2_nor2b_2 _08208_ (.A(_02630_),
    .B_N(_02711_),
    .Y(_02712_));
 sg13g2_and2_1 _08209_ (.A(_02623_),
    .B(_02712_),
    .X(_02713_));
 sg13g2_nand2_2 _08210_ (.Y(_02714_),
    .A(_02623_),
    .B(_02712_));
 sg13g2_o21ai_1 _08211_ (.B1(net3416),
    .Y(_02715_),
    .A1(net3402),
    .A2(\cpu.PC[9] ));
 sg13g2_a21oi_1 _08212_ (.A1(net3402),
    .A2(_02710_),
    .Y(_02716_),
    .B1(_02715_));
 sg13g2_nor3_2 _08213_ (.A(_02628_),
    .B(_02709_),
    .C(_02716_),
    .Y(_02717_));
 sg13g2_nand2_1 _08214_ (.Y(_02718_),
    .A(\bsq[22] ),
    .B(net3929));
 sg13g2_o21ai_1 _08215_ (.B1(_02718_),
    .Y(uio_out[7]),
    .A1(net3929),
    .A2(_02717_));
 sg13g2_o21ai_1 _08216_ (.B1(net3729),
    .Y(_02719_),
    .A1(net3734),
    .A2(_02717_));
 sg13g2_a21oi_1 _08217_ (.A1(net3734),
    .A2(uio_out[7]),
    .Y(_02720_),
    .B1(_02719_));
 sg13g2_a221oi_1 _08218_ (.B2(_01547_),
    .C1(_02720_),
    .B1(net3885),
    .A1(_01548_),
    .Y(_01308_),
    .A2(net3893));
 sg13g2_o21ai_1 _08219_ (.B1(_02119_),
    .Y(_02721_),
    .A1(_01808_),
    .A2(_02104_));
 sg13g2_nand2b_1 _08220_ (.Y(_02722_),
    .B(_02721_),
    .A_N(_02120_));
 sg13g2_mux2_2 _08221_ (.A0(\cpu.PCreg0[16] ),
    .A1(\cpu.PCreg1[16] ),
    .S(net3629),
    .X(\cpu.PC[16] ));
 sg13g2_o21ai_1 _08222_ (.B1(_02622_),
    .Y(_02723_),
    .A1(net3401),
    .A2(\cpu.PC[16] ));
 sg13g2_a21oi_1 _08223_ (.A1(net3401),
    .A2(_02722_),
    .Y(_02724_),
    .B1(_02723_));
 sg13g2_nand3_1 _08224_ (.B(_01999_),
    .C(_02015_),
    .A(_01856_),
    .Y(_02725_));
 sg13g2_nand2b_1 _08225_ (.Y(_02726_),
    .B(_02725_),
    .A_N(_02016_));
 sg13g2_mux2_2 _08226_ (.A0(\cpu.PCreg0[8] ),
    .A1(\cpu.PCreg1[8] ),
    .S(net3635),
    .X(\cpu.PC[8] ));
 sg13g2_o21ai_1 _08227_ (.B1(net3416),
    .Y(_02727_),
    .A1(net3402),
    .A2(\cpu.PC[8] ));
 sg13g2_a21oi_1 _08228_ (.A1(net3402),
    .A2(_02726_),
    .Y(_02728_),
    .B1(_02727_));
 sg13g2_mux2_1 _08229_ (.A0(_00127_),
    .A1(_00191_),
    .S(net3476),
    .X(_02729_));
 sg13g2_a21oi_1 _08230_ (.A1(net3648),
    .A2(_01692_),
    .Y(_02730_),
    .B1(net3517));
 sg13g2_o21ai_1 _08231_ (.B1(_02730_),
    .Y(_02731_),
    .A1(_00319_),
    .A2(net3511));
 sg13g2_a21oi_1 _08232_ (.A1(net3517),
    .A2(_02729_),
    .Y(_02732_),
    .B1(net3470));
 sg13g2_a21oi_1 _08233_ (.A1(_01694_),
    .A2(net3476),
    .Y(_02733_),
    .B1(net3535));
 sg13g2_o21ai_1 _08234_ (.B1(_02733_),
    .Y(_02734_),
    .A1(_00511_),
    .A2(net3476));
 sg13g2_mux2_1 _08235_ (.A0(_00159_),
    .A1(_00287_),
    .S(net3489),
    .X(_02735_));
 sg13g2_a21oi_1 _08236_ (.A1(net3538),
    .A2(_02735_),
    .Y(_02736_),
    .B1(net3465));
 sg13g2_a221oi_1 _08237_ (.B2(_02736_),
    .C1(net3461),
    .B1(_02734_),
    .A1(_02731_),
    .Y(_02737_),
    .A2(_02732_));
 sg13g2_mux4_1 _08238_ (.S0(net3477),
    .A0(_00223_),
    .A1(_00093_),
    .A2(_00383_),
    .A3(_00255_),
    .S1(net3530),
    .X(_02738_));
 sg13g2_nor2_1 _08239_ (.A(_00061_),
    .B(net3477),
    .Y(_02739_));
 sg13g2_o21ai_1 _08240_ (.B1(net3530),
    .Y(_02740_),
    .A1(net3647),
    .A2(_00351_));
 sg13g2_o21ai_1 _08241_ (.B1(net3517),
    .Y(_02741_),
    .A1(_00479_),
    .A2(net3477));
 sg13g2_o21ai_1 _08242_ (.B1(_02741_),
    .Y(_02742_),
    .A1(_02739_),
    .A2(_02740_));
 sg13g2_a221oi_1 _08243_ (.B2(net3426),
    .C1(_02737_),
    .B1(_02742_),
    .A1(net3430),
    .Y(_02743_),
    .A2(_02738_));
 sg13g2_nand2b_1 _08244_ (.Y(_02744_),
    .B(net3511),
    .A_N(_00151_));
 sg13g2_a21oi_1 _08245_ (.A1(_01652_),
    .A2(net3503),
    .Y(_02745_),
    .B1(net3547));
 sg13g2_mux2_1 _08246_ (.A0(_00471_),
    .A1(_00343_),
    .S(net3480),
    .X(_02746_));
 sg13g2_a221oi_1 _08247_ (.B2(net3532),
    .C1(net3472),
    .B1(_02746_),
    .A1(_02744_),
    .Y(_02747_),
    .A2(_02745_));
 sg13g2_mux2_1 _08248_ (.A0(_00535_),
    .A1(_00439_),
    .S(net3480),
    .X(_02748_));
 sg13g2_nand2_1 _08249_ (.Y(_02749_),
    .A(_01656_),
    .B(net3649));
 sg13g2_a21oi_1 _08250_ (.A1(_01657_),
    .A2(net3503),
    .Y(_02750_),
    .B1(net3518));
 sg13g2_a221oi_1 _08251_ (.B2(_02750_),
    .C1(net3467),
    .B1(_02749_),
    .A1(net3518),
    .Y(_02751_),
    .A2(_02748_));
 sg13g2_or3_1 _08252_ (.A(net3462),
    .B(_02747_),
    .C(_02751_),
    .X(_02752_));
 sg13g2_mux4_1 _08253_ (.S0(net3482),
    .A0(_00247_),
    .A1(_00117_),
    .A2(_00407_),
    .A3(_00279_),
    .S1(net3533),
    .X(_02753_));
 sg13g2_nor2_1 _08254_ (.A(_00085_),
    .B(net3481),
    .Y(_02754_));
 sg13g2_o21ai_1 _08255_ (.B1(net3532),
    .Y(_02755_),
    .A1(_00375_),
    .A2(net3646));
 sg13g2_o21ai_1 _08256_ (.B1(net3518),
    .Y(_02756_),
    .A1(_00503_),
    .A2(net3480));
 sg13g2_o21ai_1 _08257_ (.B1(_02756_),
    .Y(_02757_),
    .A1(_02754_),
    .A2(_02755_));
 sg13g2_a22oi_1 _08258_ (.Y(_02758_),
    .B1(_02757_),
    .B2(net3429),
    .A2(_02753_),
    .A1(net3431));
 sg13g2_and2_2 _08259_ (.A(_02752_),
    .B(_02758_),
    .X(_02759_));
 sg13g2_nand2b_1 _08260_ (.Y(_02760_),
    .B(net3515),
    .A_N(_00143_));
 sg13g2_a21oi_1 _08261_ (.A1(_01605_),
    .A2(net3500),
    .Y(_02761_),
    .B1(net3549));
 sg13g2_mux2_1 _08262_ (.A0(_00463_),
    .A1(_00335_),
    .S(net3499),
    .X(_02762_));
 sg13g2_a221oi_1 _08263_ (.B2(net3549),
    .C1(net3471),
    .B1(_02762_),
    .A1(_02760_),
    .Y(_02763_),
    .A2(_02761_));
 sg13g2_mux2_1 _08264_ (.A0(_00527_),
    .A1(_00431_),
    .S(net3499),
    .X(_02764_));
 sg13g2_nand2_1 _08265_ (.Y(_02765_),
    .A(_01608_),
    .B(net3649));
 sg13g2_a21oi_1 _08266_ (.A1(_01609_),
    .A2(net3499),
    .Y(_02766_),
    .B1(net3524));
 sg13g2_a221oi_1 _08267_ (.B2(_02766_),
    .C1(net3466),
    .B1(_02765_),
    .A1(net3524),
    .Y(_02767_),
    .A2(_02764_));
 sg13g2_or3_1 _08268_ (.A(net3463),
    .B(_02763_),
    .C(_02767_),
    .X(_02768_));
 sg13g2_mux4_1 _08269_ (.S0(net3500),
    .A0(_00239_),
    .A1(_00109_),
    .A2(_00399_),
    .A3(_00271_),
    .S1(net3546),
    .X(_02769_));
 sg13g2_nand2_1 _08270_ (.Y(_02770_),
    .A(net3433),
    .B(_02769_));
 sg13g2_nor2_1 _08271_ (.A(_00077_),
    .B(net3499),
    .Y(_02771_));
 sg13g2_o21ai_1 _08272_ (.B1(net3546),
    .Y(_02772_),
    .A1(_00367_),
    .A2(net3649));
 sg13g2_nand2_1 _08273_ (.Y(_02773_),
    .A(_00495_),
    .B(net3524));
 sg13g2_o21ai_1 _08274_ (.B1(_02773_),
    .Y(_02774_),
    .A1(_02771_),
    .A2(_02772_));
 sg13g2_nand2_1 _08275_ (.Y(_02775_),
    .A(net3427),
    .B(_02774_));
 sg13g2_nand4_1 _08276_ (.B(_02768_),
    .C(_02770_),
    .A(_02483_),
    .Y(_02776_),
    .D(_02775_));
 sg13g2_nor2_1 _08277_ (.A(net3231),
    .B(_02776_),
    .Y(_02777_));
 sg13g2_a21oi_2 _08278_ (.B1(_02777_),
    .Y(_02778_),
    .A2(net3329),
    .A1(net3231));
 sg13g2_nor2_1 _08279_ (.A(net3130),
    .B(_02778_),
    .Y(_02779_));
 sg13g2_a21oi_2 _08280_ (.B1(_02779_),
    .Y(_02780_),
    .A2(_02743_),
    .A1(net3130));
 sg13g2_nor2b_1 _08281_ (.A(_02780_),
    .B_N(net3728),
    .Y(_02781_));
 sg13g2_a21oi_1 _08282_ (.A1(_01720_),
    .A2(net3490),
    .Y(_02782_),
    .B1(net3540));
 sg13g2_o21ai_1 _08283_ (.B1(_02782_),
    .Y(_02783_),
    .A1(_00135_),
    .A2(net3490));
 sg13g2_mux2_1 _08284_ (.A0(_00455_),
    .A1(_00327_),
    .S(net3490),
    .X(_02784_));
 sg13g2_a21oi_1 _08285_ (.A1(net3540),
    .A2(_02784_),
    .Y(_02785_),
    .B1(net3469));
 sg13g2_a21oi_1 _08286_ (.A1(_01721_),
    .A2(net3490),
    .Y(_02786_),
    .B1(net3540));
 sg13g2_o21ai_1 _08287_ (.B1(_02786_),
    .Y(_02787_),
    .A1(_00519_),
    .A2(net3490));
 sg13g2_mux2_1 _08288_ (.A0(_00167_),
    .A1(_00295_),
    .S(net3490),
    .X(_02788_));
 sg13g2_a21oi_1 _08289_ (.A1(net3540),
    .A2(_02788_),
    .Y(_02789_),
    .B1(net3464));
 sg13g2_a221oi_1 _08290_ (.B2(_02789_),
    .C1(net3460),
    .B1(_02787_),
    .A1(_02783_),
    .Y(_02790_),
    .A2(_02785_));
 sg13g2_mux4_1 _08291_ (.S0(net3497),
    .A0(_00231_),
    .A1(_00101_),
    .A2(_00391_),
    .A3(_00263_),
    .S1(net3544),
    .X(_02791_));
 sg13g2_nor2_1 _08292_ (.A(_00069_),
    .B(net3497),
    .Y(_02792_));
 sg13g2_o21ai_1 _08293_ (.B1(net3544),
    .Y(_02793_),
    .A1(net3648),
    .A2(_00359_));
 sg13g2_o21ai_1 _08294_ (.B1(net3522),
    .Y(_02794_),
    .A1(_00487_),
    .A2(net3497));
 sg13g2_o21ai_1 _08295_ (.B1(_02794_),
    .Y(_02795_),
    .A1(_02792_),
    .A2(_02793_));
 sg13g2_a221oi_1 _08296_ (.B2(net3428),
    .C1(_02790_),
    .B1(_02795_),
    .A1(net3434),
    .Y(_02796_),
    .A2(_02791_));
 sg13g2_nor2b_1 _08297_ (.A(net3140),
    .B_N(_02796_),
    .Y(_02797_));
 sg13g2_a21oi_2 _08298_ (.B1(_02797_),
    .Y(_02798_),
    .A2(net3329),
    .A1(net3135));
 sg13g2_nor2_1 _08299_ (.A(net3456),
    .B(_02778_),
    .Y(_02799_));
 sg13g2_a21oi_1 _08300_ (.A1(net3723),
    .A2(net3329),
    .Y(_02800_),
    .B1(_02799_));
 sg13g2_o21ai_1 _08301_ (.B1(_02800_),
    .Y(_02801_),
    .A1(net3725),
    .A2(_02798_));
 sg13g2_nor4_2 _08302_ (.A(_02724_),
    .B(_02728_),
    .C(_02781_),
    .Y(_02802_),
    .D(_02801_));
 sg13g2_nand2_1 _08303_ (.Y(_02803_),
    .A(\bsq[21] ),
    .B(net3929));
 sg13g2_o21ai_1 _08304_ (.B1(_02803_),
    .Y(uio_out[6]),
    .A1(net3929),
    .A2(_02802_));
 sg13g2_o21ai_1 _08305_ (.B1(net3729),
    .Y(_02804_),
    .A1(net3734),
    .A2(_02802_));
 sg13g2_a21oi_1 _08306_ (.A1(net3734),
    .A2(uio_out[6]),
    .Y(_02805_),
    .B1(_02804_));
 sg13g2_a221oi_1 _08307_ (.B2(_01548_),
    .C1(_02805_),
    .B1(net3885),
    .A1(_01549_),
    .Y(_01307_),
    .A2(net3892));
 sg13g2_nor2_1 _08308_ (.A(_02408_),
    .B(_02714_),
    .Y(_02806_));
 sg13g2_xor2_1 _08309_ (.B(_02105_),
    .A(_02103_),
    .X(_02807_));
 sg13g2_mux2_2 _08310_ (.A0(\cpu.PCreg0[15] ),
    .A1(\cpu.PCreg1[15] ),
    .S(net3629),
    .X(\cpu.PC[15] ));
 sg13g2_o21ai_1 _08311_ (.B1(_02622_),
    .Y(_02808_),
    .A1(net3401),
    .A2(\cpu.PC[15] ));
 sg13g2_a21oi_1 _08312_ (.A1(net3401),
    .A2(_02807_),
    .Y(_02809_),
    .B1(_02808_));
 sg13g2_nor2_1 _08313_ (.A(_00128_),
    .B(net3497),
    .Y(_02810_));
 sg13g2_o21ai_1 _08314_ (.B1(net3522),
    .Y(_02811_),
    .A1(_00192_),
    .A2(net3513));
 sg13g2_mux2_1 _08315_ (.A0(_00448_),
    .A1(_00320_),
    .S(net3487),
    .X(_02812_));
 sg13g2_o21ai_1 _08316_ (.B1(net3468),
    .Y(_02813_),
    .A1(_02810_),
    .A2(_02811_));
 sg13g2_a21oi_1 _08317_ (.A1(net3544),
    .A2(_02812_),
    .Y(_02814_),
    .B1(_02813_));
 sg13g2_nor2_1 _08318_ (.A(_00512_),
    .B(net3488),
    .Y(_02815_));
 sg13g2_o21ai_1 _08319_ (.B1(net3521),
    .Y(_02816_),
    .A1(_00416_),
    .A2(net3512));
 sg13g2_mux2_1 _08320_ (.A0(_00160_),
    .A1(_00288_),
    .S(net3488),
    .X(_02817_));
 sg13g2_o21ai_1 _08321_ (.B1(net3470),
    .Y(_02818_),
    .A1(_02815_),
    .A2(_02816_));
 sg13g2_a21oi_1 _08322_ (.A1(net3538),
    .A2(_02817_),
    .Y(_02819_),
    .B1(_02818_));
 sg13g2_nor3_1 _08323_ (.A(net3463),
    .B(_02814_),
    .C(_02819_),
    .Y(_02820_));
 sg13g2_mux4_1 _08324_ (.S0(net3487),
    .A0(_00224_),
    .A1(_00094_),
    .A2(_00384_),
    .A3(_00256_),
    .S1(net3538),
    .X(_02821_));
 sg13g2_nor2_1 _08325_ (.A(_00062_),
    .B(net3487),
    .Y(_02822_));
 sg13g2_o21ai_1 _08326_ (.B1(net3538),
    .Y(_02823_),
    .A1(net3648),
    .A2(_00352_));
 sg13g2_o21ai_1 _08327_ (.B1(net3521),
    .Y(_02824_),
    .A1(_00480_),
    .A2(net3487));
 sg13g2_o21ai_1 _08328_ (.B1(_02824_),
    .Y(_02825_),
    .A1(_02822_),
    .A2(_02823_));
 sg13g2_a221oi_1 _08329_ (.B2(net3428),
    .C1(_02820_),
    .B1(_02825_),
    .A1(net3432),
    .Y(_02826_),
    .A2(_02821_));
 sg13g2_nand2b_1 _08330_ (.Y(_02827_),
    .B(net3514),
    .A_N(_00152_));
 sg13g2_a21oi_1 _08331_ (.A1(_01658_),
    .A2(net3509),
    .Y(_02828_),
    .B1(net3551));
 sg13g2_mux2_1 _08332_ (.A0(_00472_),
    .A1(_00344_),
    .S(net3509),
    .X(_02829_));
 sg13g2_a221oi_1 _08333_ (.B2(net3551),
    .C1(net3473),
    .B1(_02829_),
    .A1(_02827_),
    .Y(_02830_),
    .A2(_02828_));
 sg13g2_mux2_1 _08334_ (.A0(_00536_),
    .A1(_00440_),
    .S(net3507),
    .X(_02831_));
 sg13g2_nand2_1 _08335_ (.Y(_02832_),
    .A(_01662_),
    .B(net3650));
 sg13g2_a21oi_1 _08336_ (.A1(_01663_),
    .A2(net3507),
    .Y(_02833_),
    .B1(net3526));
 sg13g2_a221oi_1 _08337_ (.B2(_02833_),
    .C1(net3466),
    .B1(_02832_),
    .A1(net3526),
    .Y(_02834_),
    .A2(_02831_));
 sg13g2_or3_2 _08338_ (.A(net3462),
    .B(_02830_),
    .C(_02834_),
    .X(_02835_));
 sg13g2_mux4_1 _08339_ (.S0(net3502),
    .A0(_00248_),
    .A1(_00118_),
    .A2(_00408_),
    .A3(_00280_),
    .S1(net3547),
    .X(_02836_));
 sg13g2_nor2_1 _08340_ (.A(_00086_),
    .B(net3502),
    .Y(_02837_));
 sg13g2_o21ai_1 _08341_ (.B1(net3548),
    .Y(_02838_),
    .A1(_00376_),
    .A2(net3649));
 sg13g2_o21ai_1 _08342_ (.B1(net3525),
    .Y(_02839_),
    .A1(_00504_),
    .A2(net3502));
 sg13g2_o21ai_1 _08343_ (.B1(_02839_),
    .Y(_02840_),
    .A1(_02837_),
    .A2(_02838_));
 sg13g2_a22oi_1 _08344_ (.Y(_02841_),
    .B1(_02840_),
    .B2(net3427),
    .A2(_02836_),
    .A1(net3433));
 sg13g2_and2_2 _08345_ (.A(_02835_),
    .B(_02841_),
    .X(_02842_));
 sg13g2_nand2b_1 _08346_ (.Y(_02843_),
    .B(net3511),
    .A_N(_00144_));
 sg13g2_a21oi_1 _08347_ (.A1(_01610_),
    .A2(net3486),
    .Y(_02844_),
    .B1(net3536));
 sg13g2_mux2_1 _08348_ (.A0(_00464_),
    .A1(_00336_),
    .S(net3486),
    .X(_02845_));
 sg13g2_a221oi_1 _08349_ (.B2(net3536),
    .C1(net3470),
    .B1(_02845_),
    .A1(_02843_),
    .Y(_02846_),
    .A2(_02844_));
 sg13g2_mux2_1 _08350_ (.A0(_00528_),
    .A1(_00432_),
    .S(net3484),
    .X(_02847_));
 sg13g2_nand2b_1 _08351_ (.Y(_02848_),
    .B(net3648),
    .A_N(_00176_));
 sg13g2_a21oi_1 _08352_ (.A1(_01615_),
    .A2(net3486),
    .Y(_02849_),
    .B1(net3521));
 sg13g2_a221oi_1 _08353_ (.B2(_02849_),
    .C1(net3465),
    .B1(_02848_),
    .A1(net3521),
    .Y(_02850_),
    .A2(_02847_));
 sg13g2_or3_1 _08354_ (.A(net3461),
    .B(_02846_),
    .C(_02850_),
    .X(_02851_));
 sg13g2_mux4_1 _08355_ (.S0(net3477),
    .A0(_00240_),
    .A1(_00110_),
    .A2(_00400_),
    .A3(_00272_),
    .S1(net3530),
    .X(_02852_));
 sg13g2_nand2_1 _08356_ (.Y(_02853_),
    .A(net3430),
    .B(_02852_));
 sg13g2_nor2_1 _08357_ (.A(_00078_),
    .B(net3477),
    .Y(_02854_));
 sg13g2_o21ai_1 _08358_ (.B1(net3530),
    .Y(_02855_),
    .A1(_00368_),
    .A2(net3647));
 sg13g2_nand2_1 _08359_ (.Y(_02856_),
    .A(_00496_),
    .B(net3517));
 sg13g2_o21ai_1 _08360_ (.B1(_02856_),
    .Y(_02857_),
    .A1(_02854_),
    .A2(_02855_));
 sg13g2_nand2_1 _08361_ (.Y(_02858_),
    .A(net3426),
    .B(_02857_));
 sg13g2_nand4_1 _08362_ (.B(_02851_),
    .C(_02853_),
    .A(_02483_),
    .Y(_02859_),
    .D(_02858_));
 sg13g2_nor2_1 _08363_ (.A(net3231),
    .B(_02859_),
    .Y(_02860_));
 sg13g2_a21oi_2 _08364_ (.B1(_02860_),
    .Y(_02861_),
    .A2(net3328),
    .A1(net3231));
 sg13g2_nor2_1 _08365_ (.A(net3131),
    .B(_02861_),
    .Y(_02862_));
 sg13g2_a21oi_2 _08366_ (.B1(_02862_),
    .Y(_02863_),
    .A2(_02826_),
    .A1(net3131));
 sg13g2_nor2b_1 _08367_ (.A(_02863_),
    .B_N(net3728),
    .Y(_02864_));
 sg13g2_a21oi_1 _08368_ (.A1(_01576_),
    .A2(net3493),
    .Y(_02865_),
    .B1(net3545));
 sg13g2_o21ai_1 _08369_ (.B1(_02865_),
    .Y(_02866_),
    .A1(_00136_),
    .A2(net3493));
 sg13g2_mux2_1 _08370_ (.A0(_00456_),
    .A1(_00328_),
    .S(net3493),
    .X(_02867_));
 sg13g2_a21oi_1 _08371_ (.A1(net3541),
    .A2(_02867_),
    .Y(_02868_),
    .B1(net3469));
 sg13g2_o21ai_1 _08372_ (.B1(net3522),
    .Y(_02869_),
    .A1(_00424_),
    .A2(net3513));
 sg13g2_a21o_1 _08373_ (.A2(net3513),
    .A1(_01579_),
    .B1(_02869_),
    .X(_02870_));
 sg13g2_mux2_1 _08374_ (.A0(_00168_),
    .A1(_00296_),
    .S(net3493),
    .X(_02871_));
 sg13g2_a21oi_1 _08375_ (.A1(net3541),
    .A2(_02871_),
    .Y(_02872_),
    .B1(net3464));
 sg13g2_a221oi_1 _08376_ (.B2(_02872_),
    .C1(net3460),
    .B1(_02870_),
    .A1(_02866_),
    .Y(_02873_),
    .A2(_02868_));
 sg13g2_mux4_1 _08377_ (.S0(net3493),
    .A0(_00232_),
    .A1(_00102_),
    .A2(_00392_),
    .A3(_00264_),
    .S1(net3541),
    .X(_02874_));
 sg13g2_nor2_1 _08378_ (.A(_00070_),
    .B(net3493),
    .Y(_02875_));
 sg13g2_o21ai_1 _08379_ (.B1(net3541),
    .Y(_02876_),
    .A1(_00360_),
    .A2(net3652));
 sg13g2_o21ai_1 _08380_ (.B1(net3522),
    .Y(_02877_),
    .A1(_00488_),
    .A2(net3493));
 sg13g2_o21ai_1 _08381_ (.B1(_02877_),
    .Y(_02878_),
    .A1(_02875_),
    .A2(_02876_));
 sg13g2_a221oi_1 _08382_ (.B2(net3428),
    .C1(_02873_),
    .B1(_02878_),
    .A1(net3432),
    .Y(_02879_),
    .A2(_02874_));
 sg13g2_nor2b_1 _08383_ (.A(net3135),
    .B_N(_02879_),
    .Y(_02880_));
 sg13g2_a21oi_2 _08384_ (.B1(_02880_),
    .Y(_02881_),
    .A2(net3328),
    .A1(net3135));
 sg13g2_nor2_1 _08385_ (.A(net3725),
    .B(_02881_),
    .Y(_02882_));
 sg13g2_a21oi_1 _08386_ (.A1(net3723),
    .A2(net3328),
    .Y(_02883_),
    .B1(net3416));
 sg13g2_o21ai_1 _08387_ (.B1(_02883_),
    .Y(_02884_),
    .A1(net3456),
    .A2(_02861_));
 sg13g2_nor4_2 _08388_ (.A(_02809_),
    .B(_02864_),
    .C(_02882_),
    .Y(_02885_),
    .D(_02884_));
 sg13g2_nor2_2 _08389_ (.A(_02806_),
    .B(_02885_),
    .Y(_02886_));
 sg13g2_mux2_2 _08390_ (.A0(_02886_),
    .A1(\bsq[20] ),
    .S(net3930),
    .X(uio_out[5]));
 sg13g2_nor2_1 _08391_ (.A(net3735),
    .B(_02886_),
    .Y(_02887_));
 sg13g2_o21ai_1 _08392_ (.B1(net3729),
    .Y(_02888_),
    .A1(net3900),
    .A2(uio_out[5]));
 sg13g2_a21oi_1 _08393_ (.A1(\jtag0.bssh[21] ),
    .A2(net3927),
    .Y(_02889_),
    .B1(net3892));
 sg13g2_o21ai_1 _08394_ (.B1(_02889_),
    .Y(_02890_),
    .A1(_02887_),
    .A2(_02888_));
 sg13g2_o21ai_1 _08395_ (.B1(_02890_),
    .Y(_02891_),
    .A1(\jtag0.bssh[20] ),
    .A2(_02586_));
 sg13g2_inv_1 _08396_ (.Y(_01306_),
    .A(_02891_));
 sg13g2_xnor2_1 _08397_ (.Y(_02892_),
    .A(_02101_),
    .B(_02102_));
 sg13g2_mux2_2 _08398_ (.A0(\cpu.PCreg0[14] ),
    .A1(\cpu.PCreg1[14] ),
    .S(net3629),
    .X(\cpu.PC[14] ));
 sg13g2_a21oi_1 _08399_ (.A1(net3405),
    .A2(_02892_),
    .Y(_02893_),
    .B1(_02623_));
 sg13g2_o21ai_1 _08400_ (.B1(_02893_),
    .Y(_02894_),
    .A1(net3402),
    .A2(\cpu.PC[14] ));
 sg13g2_nor2_1 _08401_ (.A(_00129_),
    .B(net3487),
    .Y(_02895_));
 sg13g2_o21ai_1 _08402_ (.B1(net3523),
    .Y(_02896_),
    .A1(_00193_),
    .A2(net3512));
 sg13g2_mux2_1 _08403_ (.A0(_00449_),
    .A1(_00321_),
    .S(net3487),
    .X(_02897_));
 sg13g2_o21ai_1 _08404_ (.B1(net3465),
    .Y(_02898_),
    .A1(_02895_),
    .A2(_02896_));
 sg13g2_a21oi_1 _08405_ (.A1(net3539),
    .A2(_02897_),
    .Y(_02899_),
    .B1(_02898_));
 sg13g2_nor2_1 _08406_ (.A(_00513_),
    .B(net3485),
    .Y(_02900_));
 sg13g2_o21ai_1 _08407_ (.B1(net3521),
    .Y(_02901_),
    .A1(_00417_),
    .A2(net3512));
 sg13g2_mux2_1 _08408_ (.A0(_00161_),
    .A1(_00289_),
    .S(net3485),
    .X(_02902_));
 sg13g2_o21ai_1 _08409_ (.B1(net3469),
    .Y(_02903_),
    .A1(_02900_),
    .A2(_02901_));
 sg13g2_a21oi_1 _08410_ (.A1(net3539),
    .A2(_02902_),
    .Y(_02904_),
    .B1(_02903_));
 sg13g2_nor3_1 _08411_ (.A(net3463),
    .B(_02899_),
    .C(_02904_),
    .Y(_02905_));
 sg13g2_mux4_1 _08412_ (.S0(net3489),
    .A0(_00225_),
    .A1(_00095_),
    .A2(_00385_),
    .A3(_00257_),
    .S1(net3538),
    .X(_02906_));
 sg13g2_nor2_1 _08413_ (.A(_00063_),
    .B(net3488),
    .Y(_02907_));
 sg13g2_o21ai_1 _08414_ (.B1(net3538),
    .Y(_02908_),
    .A1(net3648),
    .A2(_00353_));
 sg13g2_o21ai_1 _08415_ (.B1(net3523),
    .Y(_02909_),
    .A1(_00481_),
    .A2(net3488));
 sg13g2_o21ai_1 _08416_ (.B1(_02909_),
    .Y(_02910_),
    .A1(_02907_),
    .A2(_02908_));
 sg13g2_a221oi_1 _08417_ (.B2(net3428),
    .C1(_02905_),
    .B1(_02910_),
    .A1(net3432),
    .Y(_02911_),
    .A2(_02906_));
 sg13g2_nand2b_1 _08418_ (.Y(_02912_),
    .B(net3516),
    .A_N(_00153_));
 sg13g2_a21oi_1 _08419_ (.A1(_01665_),
    .A2(net3481),
    .Y(_02913_),
    .B1(net3531));
 sg13g2_mux2_1 _08420_ (.A0(_00473_),
    .A1(_00345_),
    .S(net3478),
    .X(_02914_));
 sg13g2_a221oi_1 _08421_ (.B2(net3531),
    .C1(net3472),
    .B1(_02914_),
    .A1(_02912_),
    .Y(_02915_),
    .A2(_02913_));
 sg13g2_mux2_1 _08422_ (.A0(_00537_),
    .A1(_00441_),
    .S(net3478),
    .X(_02916_));
 sg13g2_nand2_1 _08423_ (.Y(_02917_),
    .A(_01669_),
    .B(net3645));
 sg13g2_a21oi_1 _08424_ (.A1(_01670_),
    .A2(net3478),
    .Y(_02918_),
    .B1(net3519));
 sg13g2_a221oi_1 _08425_ (.B2(_02918_),
    .C1(net3467),
    .B1(_02917_),
    .A1(net3519),
    .Y(_02919_),
    .A2(_02916_));
 sg13g2_or3_2 _08426_ (.A(net3462),
    .B(_02915_),
    .C(_02919_),
    .X(_02920_));
 sg13g2_mux4_1 _08427_ (.S0(net3478),
    .A0(_00249_),
    .A1(_00119_),
    .A2(_00409_),
    .A3(_00281_),
    .S1(net3531),
    .X(_02921_));
 sg13g2_nor2_1 _08428_ (.A(_00087_),
    .B(net3478),
    .Y(_02922_));
 sg13g2_o21ai_1 _08429_ (.B1(net3531),
    .Y(_02923_),
    .A1(_00377_),
    .A2(net3646));
 sg13g2_o21ai_1 _08430_ (.B1(net3519),
    .Y(_02924_),
    .A1(_00505_),
    .A2(net3478));
 sg13g2_o21ai_1 _08431_ (.B1(_02924_),
    .Y(_02925_),
    .A1(_02922_),
    .A2(_02923_));
 sg13g2_a22oi_1 _08432_ (.Y(_02926_),
    .B1(_02925_),
    .B2(net3426),
    .A2(_02921_),
    .A1(net3430));
 sg13g2_and2_2 _08433_ (.A(_02920_),
    .B(_02926_),
    .X(_02927_));
 sg13g2_nand2_2 _08434_ (.Y(_02928_),
    .A(_02920_),
    .B(_02926_));
 sg13g2_nand2b_1 _08435_ (.Y(_02929_),
    .B(net3511),
    .A_N(_00145_));
 sg13g2_a21oi_1 _08436_ (.A1(_01616_),
    .A2(net3474),
    .Y(_02930_),
    .B1(net3529));
 sg13g2_mux2_1 _08437_ (.A0(_00465_),
    .A1(_00337_),
    .S(net3475),
    .X(_02931_));
 sg13g2_a221oi_1 _08438_ (.B2(net3529),
    .C1(net3470),
    .B1(_02931_),
    .A1(_02929_),
    .Y(_02932_),
    .A2(_02930_));
 sg13g2_mux2_1 _08439_ (.A0(_00529_),
    .A1(_00433_),
    .S(net3474),
    .X(_02933_));
 sg13g2_nand2b_1 _08440_ (.Y(_02934_),
    .B(net3647),
    .A_N(_00177_));
 sg13g2_a21oi_1 _08441_ (.A1(_01621_),
    .A2(net3474),
    .Y(_02935_),
    .B1(net3517));
 sg13g2_a221oi_1 _08442_ (.B2(_02935_),
    .C1(net3465),
    .B1(_02934_),
    .A1(net3517),
    .Y(_02936_),
    .A2(_02933_));
 sg13g2_or3_1 _08443_ (.A(net3461),
    .B(_02932_),
    .C(_02936_),
    .X(_02937_));
 sg13g2_mux4_1 _08444_ (.S0(net3477),
    .A0(_00241_),
    .A1(_00111_),
    .A2(_00401_),
    .A3(_00273_),
    .S1(net3530),
    .X(_02938_));
 sg13g2_nand2_1 _08445_ (.Y(_02939_),
    .A(net3430),
    .B(_02938_));
 sg13g2_nor2_1 _08446_ (.A(_00079_),
    .B(net3475),
    .Y(_02940_));
 sg13g2_o21ai_1 _08447_ (.B1(net3530),
    .Y(_02941_),
    .A1(_00369_),
    .A2(net3647));
 sg13g2_nand2_1 _08448_ (.Y(_02942_),
    .A(_00497_),
    .B(net3517));
 sg13g2_o21ai_1 _08449_ (.B1(_02942_),
    .Y(_02943_),
    .A1(_02940_),
    .A2(_02941_));
 sg13g2_nand2_1 _08450_ (.Y(_02944_),
    .A(net3426),
    .B(_02943_));
 sg13g2_nand4_1 _08451_ (.B(_02937_),
    .C(_02939_),
    .A(_02483_),
    .Y(_02945_),
    .D(_02944_));
 sg13g2_nor2_1 _08452_ (.A(net3232),
    .B(_02945_),
    .Y(_02946_));
 sg13g2_a21oi_2 _08453_ (.B1(_02946_),
    .Y(_02947_),
    .A2(_02927_),
    .A1(net3231));
 sg13g2_nor2_1 _08454_ (.A(net3130),
    .B(_02947_),
    .Y(_02948_));
 sg13g2_a21oi_2 _08455_ (.B1(_02948_),
    .Y(_02949_),
    .A2(_02911_),
    .A1(net3130));
 sg13g2_nor2b_1 _08456_ (.A(_02949_),
    .B_N(net3728),
    .Y(_02950_));
 sg13g2_a21oi_1 _08457_ (.A1(_01580_),
    .A2(net3484),
    .Y(_02951_),
    .B1(net3536));
 sg13g2_o21ai_1 _08458_ (.B1(_02951_),
    .Y(_02952_),
    .A1(_00137_),
    .A2(net3484));
 sg13g2_mux2_1 _08459_ (.A0(_00457_),
    .A1(_00329_),
    .S(net3484),
    .X(_02953_));
 sg13g2_a21oi_1 _08460_ (.A1(net3536),
    .A2(_02953_),
    .Y(_02954_),
    .B1(net3470));
 sg13g2_a21oi_1 _08461_ (.A1(_01581_),
    .A2(net3484),
    .Y(_02955_),
    .B1(net3536));
 sg13g2_o21ai_1 _08462_ (.B1(_02955_),
    .Y(_02956_),
    .A1(_00521_),
    .A2(net3484));
 sg13g2_mux2_1 _08463_ (.A0(_00169_),
    .A1(_00297_),
    .S(net3484),
    .X(_02957_));
 sg13g2_a21oi_1 _08464_ (.A1(net3536),
    .A2(_02957_),
    .Y(_02958_),
    .B1(net3465));
 sg13g2_a221oi_1 _08465_ (.B2(_02958_),
    .C1(net3461),
    .B1(_02956_),
    .A1(_02952_),
    .Y(_02959_),
    .A2(_02954_));
 sg13g2_mux4_1 _08466_ (.S0(net3477),
    .A0(_00233_),
    .A1(_00103_),
    .A2(_00393_),
    .A3(_00265_),
    .S1(net3530),
    .X(_02960_));
 sg13g2_nor2_1 _08467_ (.A(_00071_),
    .B(net3475),
    .Y(_02961_));
 sg13g2_o21ai_1 _08468_ (.B1(net3529),
    .Y(_02962_),
    .A1(_00361_),
    .A2(net3647));
 sg13g2_o21ai_1 _08469_ (.B1(net3520),
    .Y(_02963_),
    .A1(_00489_),
    .A2(net3475));
 sg13g2_o21ai_1 _08470_ (.B1(_02963_),
    .Y(_02964_),
    .A1(_02961_),
    .A2(_02962_));
 sg13g2_a221oi_1 _08471_ (.B2(net3426),
    .C1(_02959_),
    .B1(_02964_),
    .A1(net3430),
    .Y(_02965_),
    .A2(_02960_));
 sg13g2_nand2_1 _08472_ (.Y(_02966_),
    .A(net3135),
    .B(_02928_));
 sg13g2_o21ai_1 _08473_ (.B1(_02966_),
    .Y(_02967_),
    .A1(net3135),
    .A2(_02965_));
 sg13g2_nor2_1 _08474_ (.A(net3725),
    .B(_02967_),
    .Y(_02968_));
 sg13g2_a21oi_1 _08475_ (.A1(net3723),
    .A2(_02927_),
    .Y(_02969_),
    .B1(net3416));
 sg13g2_o21ai_1 _08476_ (.B1(_02969_),
    .Y(_02970_),
    .A1(net3456),
    .A2(_02947_));
 sg13g2_nor3_1 _08477_ (.A(_02950_),
    .B(_02968_),
    .C(_02970_),
    .Y(_02971_));
 sg13g2_a22oi_1 _08478_ (.Y(_02972_),
    .B1(_02894_),
    .B2(_02971_),
    .A2(_02713_),
    .A1(net3119));
 sg13g2_mux2_2 _08479_ (.A0(_02972_),
    .A1(\bsq[19] ),
    .S(net3930),
    .X(uio_out[4]));
 sg13g2_nor2_1 _08480_ (.A(net3735),
    .B(_02972_),
    .Y(_02973_));
 sg13g2_o21ai_1 _08481_ (.B1(net3729),
    .Y(_02974_),
    .A1(net3900),
    .A2(uio_out[4]));
 sg13g2_a21oi_1 _08482_ (.A1(\jtag0.bssh[20] ),
    .A2(net3927),
    .Y(_02975_),
    .B1(net3892));
 sg13g2_o21ai_1 _08483_ (.B1(_02975_),
    .Y(_02976_),
    .A1(_02973_),
    .A2(_02974_));
 sg13g2_o21ai_1 _08484_ (.B1(_02976_),
    .Y(_02977_),
    .A1(\jtag0.bssh[19] ),
    .A2(_02586_));
 sg13g2_inv_1 _08485_ (.Y(_01305_),
    .A(_02977_));
 sg13g2_mux2_2 _08486_ (.A0(\cpu.PCreg0[13] ),
    .A1(\cpu.PCreg1[13] ),
    .S(net3629),
    .X(\cpu.PC[13] ));
 sg13g2_o21ai_1 _08487_ (.B1(_02622_),
    .Y(_02978_),
    .A1(net3401),
    .A2(\cpu.PC[13] ));
 sg13g2_a21oi_1 _08488_ (.A1(net3628),
    .A2(_02078_),
    .Y(_02979_),
    .B1(_02081_));
 sg13g2_xor2_1 _08489_ (.B(_02979_),
    .A(_02098_),
    .X(_02980_));
 sg13g2_nor2_1 _08490_ (.A(net3407),
    .B(_02980_),
    .Y(_02981_));
 sg13g2_a21oi_1 _08491_ (.A1(_01719_),
    .A2(net3492),
    .Y(_02982_),
    .B1(net3541));
 sg13g2_o21ai_1 _08492_ (.B1(_02982_),
    .Y(_02983_),
    .A1(_00130_),
    .A2(net3492));
 sg13g2_mux2_1 _08493_ (.A0(_00450_),
    .A1(_00322_),
    .S(net3492),
    .X(_02984_));
 sg13g2_a21oi_1 _08494_ (.A1(net3541),
    .A2(_02984_),
    .Y(_02985_),
    .B1(net3469));
 sg13g2_nor2_1 _08495_ (.A(_00514_),
    .B(net3497),
    .Y(_02986_));
 sg13g2_o21ai_1 _08496_ (.B1(net3522),
    .Y(_02987_),
    .A1(_00418_),
    .A2(net3513));
 sg13g2_mux2_1 _08497_ (.A0(_00162_),
    .A1(_00290_),
    .S(net3497),
    .X(_02988_));
 sg13g2_a21oi_1 _08498_ (.A1(net3544),
    .A2(_02988_),
    .Y(_02989_),
    .B1(net3468));
 sg13g2_o21ai_1 _08499_ (.B1(_02989_),
    .Y(_02990_),
    .A1(_02986_),
    .A2(_02987_));
 sg13g2_a21oi_1 _08500_ (.A1(_02983_),
    .A2(_02985_),
    .Y(_02991_),
    .B1(net3460));
 sg13g2_mux4_1 _08501_ (.S0(net3487),
    .A0(_00226_),
    .A1(_00096_),
    .A2(_00386_),
    .A3(_00258_),
    .S1(net3538),
    .X(_02992_));
 sg13g2_o21ai_1 _08502_ (.B1(net3544),
    .Y(_02993_),
    .A1(net3648),
    .A2(_00354_));
 sg13g2_a21oi_1 _08503_ (.A1(_01718_),
    .A2(net3513),
    .Y(_02994_),
    .B1(_02993_));
 sg13g2_a21oi_1 _08504_ (.A1(_00482_),
    .A2(net3522),
    .Y(_02995_),
    .B1(_02994_));
 sg13g2_o21ai_1 _08505_ (.B1(_02483_),
    .Y(_02996_),
    .A1(_02463_),
    .A2(_02995_));
 sg13g2_a221oi_1 _08506_ (.B2(net3434),
    .C1(_02996_),
    .B1(_02992_),
    .A1(_02990_),
    .Y(_02997_),
    .A2(_02991_));
 sg13g2_nand2b_1 _08507_ (.Y(_02998_),
    .B(net3515),
    .A_N(_00154_));
 sg13g2_a21oi_1 _08508_ (.A1(_01671_),
    .A2(net3501),
    .Y(_02999_),
    .B1(net3548));
 sg13g2_mux2_1 _08509_ (.A0(_00474_),
    .A1(_00346_),
    .S(net3501),
    .X(_03000_));
 sg13g2_a221oi_1 _08510_ (.B2(net3548),
    .C1(net3471),
    .B1(_03000_),
    .A1(_02998_),
    .Y(_03001_),
    .A2(_02999_));
 sg13g2_nand2b_1 _08511_ (.Y(_03002_),
    .B(net3515),
    .A_N(_00538_));
 sg13g2_a21oi_1 _08512_ (.A1(_01674_),
    .A2(net3501),
    .Y(_03003_),
    .B1(net3548));
 sg13g2_mux2_1 _08513_ (.A0(_00186_),
    .A1(_00314_),
    .S(net3501),
    .X(_03004_));
 sg13g2_a221oi_1 _08514_ (.B2(net3548),
    .C1(net3466),
    .B1(_03004_),
    .A1(_03002_),
    .Y(_03005_),
    .A2(_03003_));
 sg13g2_or3_2 _08515_ (.A(net3462),
    .B(_03001_),
    .C(_03005_),
    .X(_03006_));
 sg13g2_mux4_1 _08516_ (.S0(net3480),
    .A0(_00250_),
    .A1(_00120_),
    .A2(_00410_),
    .A3(_00282_),
    .S1(net3547),
    .X(_03007_));
 sg13g2_nand2_1 _08517_ (.Y(_03008_),
    .A(net3431),
    .B(_03007_));
 sg13g2_nand2_1 _08518_ (.Y(_03009_),
    .A(_00506_),
    .B(net3524));
 sg13g2_nor2_1 _08519_ (.A(_00088_),
    .B(net3503),
    .Y(_03010_));
 sg13g2_o21ai_1 _08520_ (.B1(net3547),
    .Y(_03011_),
    .A1(_00378_),
    .A2(net3649));
 sg13g2_o21ai_1 _08521_ (.B1(_03009_),
    .Y(_03012_),
    .A1(_03010_),
    .A2(_03011_));
 sg13g2_a21oi_2 _08522_ (.B1(net3386),
    .Y(_03013_),
    .A2(_03012_),
    .A1(net3427));
 sg13g2_and3_2 _08523_ (.X(_03014_),
    .A(_03006_),
    .B(_03008_),
    .C(_03013_));
 sg13g2_nand2b_1 _08524_ (.Y(_03015_),
    .B(net3514),
    .A_N(_00146_));
 sg13g2_a21oi_1 _08525_ (.A1(_01622_),
    .A2(net3505),
    .Y(_03016_),
    .B1(net3550));
 sg13g2_mux2_1 _08526_ (.A0(_00466_),
    .A1(_00338_),
    .S(net3505),
    .X(_03017_));
 sg13g2_a221oi_1 _08527_ (.B2(net3550),
    .C1(net3471),
    .B1(_03017_),
    .A1(_03015_),
    .Y(_03018_),
    .A2(_03016_));
 sg13g2_nor2_1 _08528_ (.A(_00530_),
    .B(net3505),
    .Y(_03019_));
 sg13g2_a21oi_1 _08529_ (.A1(_01625_),
    .A2(net3505),
    .Y(_03020_),
    .B1(_03019_));
 sg13g2_nand2_1 _08530_ (.Y(_03021_),
    .A(_01626_),
    .B(net3650));
 sg13g2_a21oi_1 _08531_ (.A1(_01627_),
    .A2(net3505),
    .Y(_03022_),
    .B1(net3527));
 sg13g2_a221oi_1 _08532_ (.B2(_03022_),
    .C1(net3466),
    .B1(_03021_),
    .A1(net3527),
    .Y(_03023_),
    .A2(_03020_));
 sg13g2_nand2b_1 _08533_ (.Y(_03024_),
    .B(_02452_),
    .A_N(_03018_));
 sg13g2_mux4_1 _08534_ (.S0(net3506),
    .A0(_00242_),
    .A1(_00112_),
    .A2(_00402_),
    .A3(_00274_),
    .S1(net3552),
    .X(_03025_));
 sg13g2_nand2_1 _08535_ (.Y(_03026_),
    .A(_00498_),
    .B(net3527));
 sg13g2_nor2_1 _08536_ (.A(_00080_),
    .B(net3505),
    .Y(_03027_));
 sg13g2_o21ai_1 _08537_ (.B1(net3550),
    .Y(_03028_),
    .A1(_00370_),
    .A2(net3650));
 sg13g2_o21ai_1 _08538_ (.B1(_03026_),
    .Y(_03029_),
    .A1(_03027_),
    .A2(_03028_));
 sg13g2_a221oi_1 _08539_ (.B2(net3427),
    .C1(net3386),
    .B1(_03029_),
    .A1(net3434),
    .Y(_03030_),
    .A2(_03025_));
 sg13g2_o21ai_1 _08540_ (.B1(_03030_),
    .Y(_03031_),
    .A1(_03023_),
    .A2(_03024_));
 sg13g2_nor2_1 _08541_ (.A(net3232),
    .B(_03031_),
    .Y(_03032_));
 sg13g2_a21oi_2 _08542_ (.B1(_03032_),
    .Y(_03033_),
    .A2(_03014_),
    .A1(net3232));
 sg13g2_nor2_1 _08543_ (.A(net3130),
    .B(_03033_),
    .Y(_03034_));
 sg13g2_a21oi_2 _08544_ (.B1(_03034_),
    .Y(_03035_),
    .A2(_02997_),
    .A1(net3131));
 sg13g2_nor2b_1 _08545_ (.A(_03035_),
    .B_N(net3728),
    .Y(_03036_));
 sg13g2_a21oi_1 _08546_ (.A1(_01582_),
    .A2(net3494),
    .Y(_03037_),
    .B1(net3542));
 sg13g2_o21ai_1 _08547_ (.B1(_03037_),
    .Y(_03038_),
    .A1(_00138_),
    .A2(net3494));
 sg13g2_mux2_1 _08548_ (.A0(_00458_),
    .A1(_00330_),
    .S(net3495),
    .X(_03039_));
 sg13g2_a21oi_1 _08549_ (.A1(net3542),
    .A2(_03039_),
    .Y(_03040_),
    .B1(net3469));
 sg13g2_a21oi_1 _08550_ (.A1(_01586_),
    .A2(net3494),
    .Y(_03041_),
    .B1(net3542));
 sg13g2_o21ai_1 _08551_ (.B1(_03041_),
    .Y(_03042_),
    .A1(_00522_),
    .A2(net3494));
 sg13g2_mux2_1 _08552_ (.A0(_00170_),
    .A1(_00298_),
    .S(net3494),
    .X(_03043_));
 sg13g2_a21oi_1 _08553_ (.A1(net3542),
    .A2(_03043_),
    .Y(_03044_),
    .B1(net3464));
 sg13g2_a221oi_1 _08554_ (.B2(_03044_),
    .C1(net3460),
    .B1(_03042_),
    .A1(_03038_),
    .Y(_03045_),
    .A2(_03040_));
 sg13g2_mux4_1 _08555_ (.S0(net3497),
    .A0(_00234_),
    .A1(_00104_),
    .A2(_00394_),
    .A3(_00266_),
    .S1(net3544),
    .X(_03046_));
 sg13g2_nand2_1 _08556_ (.Y(_03047_),
    .A(_00490_),
    .B(net3527));
 sg13g2_nor2_1 _08557_ (.A(_00072_),
    .B(net3505),
    .Y(_03048_));
 sg13g2_o21ai_1 _08558_ (.B1(net3542),
    .Y(_03049_),
    .A1(_00362_),
    .A2(net3648));
 sg13g2_o21ai_1 _08559_ (.B1(_03047_),
    .Y(_03050_),
    .A1(_03048_),
    .A2(_03049_));
 sg13g2_a221oi_1 _08560_ (.B2(net3428),
    .C1(_02482_),
    .B1(_03050_),
    .A1(net3432),
    .Y(_03051_),
    .A2(_03046_));
 sg13g2_nand2b_2 _08561_ (.Y(_03052_),
    .B(_03051_),
    .A_N(_03045_));
 sg13g2_nor2_1 _08562_ (.A(net3136),
    .B(_03052_),
    .Y(_03053_));
 sg13g2_a21oi_2 _08563_ (.B1(_03053_),
    .Y(_03054_),
    .A2(net3327),
    .A1(net3136));
 sg13g2_nor2_1 _08564_ (.A(net3725),
    .B(_03054_),
    .Y(_03055_));
 sg13g2_a21oi_1 _08565_ (.A1(net3723),
    .A2(net3327),
    .Y(_03056_),
    .B1(net3416));
 sg13g2_o21ai_1 _08566_ (.B1(_03056_),
    .Y(_03057_),
    .A1(net3456),
    .A2(_03033_));
 sg13g2_nor3_1 _08567_ (.A(_03036_),
    .B(_03055_),
    .C(_03057_),
    .Y(_03058_));
 sg13g2_o21ai_1 _08568_ (.B1(_03058_),
    .Y(_03059_),
    .A1(_02978_),
    .A2(_02981_));
 sg13g2_o21ai_1 _08569_ (.B1(_03059_),
    .Y(_03060_),
    .A1(net3128),
    .A2(_02714_));
 sg13g2_nand2_1 _08570_ (.Y(_03061_),
    .A(\bsq[18] ),
    .B(net3931));
 sg13g2_o21ai_1 _08571_ (.B1(_03061_),
    .Y(uio_out[3]),
    .A1(net3930),
    .A2(_03060_));
 sg13g2_a21oi_1 _08572_ (.A1(net3900),
    .A2(_03060_),
    .Y(_03062_),
    .B1(_02589_));
 sg13g2_o21ai_1 _08573_ (.B1(_03062_),
    .Y(_03063_),
    .A1(net3900),
    .A2(uio_out[3]));
 sg13g2_a21oi_1 _08574_ (.A1(\jtag0.bssh[19] ),
    .A2(net3928),
    .Y(_03064_),
    .B1(net3896));
 sg13g2_a22oi_1 _08575_ (.Y(_01304_),
    .B1(_03063_),
    .B2(_03064_),
    .A2(net3896),
    .A1(_01550_));
 sg13g2_nor3_1 _08576_ (.A(_02060_),
    .B(_02062_),
    .C(_02080_),
    .Y(_03065_));
 sg13g2_or2_1 _08577_ (.X(_03066_),
    .B(_03065_),
    .A(_02081_));
 sg13g2_mux2_2 _08578_ (.A0(\cpu.PCreg0[12] ),
    .A1(\cpu.PCreg1[12] ),
    .S(net3629),
    .X(\cpu.PC[12] ));
 sg13g2_o21ai_1 _08579_ (.B1(_02622_),
    .Y(_03067_),
    .A1(net3401),
    .A2(\cpu.PC[12] ));
 sg13g2_a21oi_1 _08580_ (.A1(net3403),
    .A2(_03066_),
    .Y(_03068_),
    .B1(_03067_));
 sg13g2_a21oi_1 _08581_ (.A1(_01716_),
    .A2(net3474),
    .Y(_03069_),
    .B1(net3529));
 sg13g2_o21ai_1 _08582_ (.B1(_03069_),
    .Y(_03070_),
    .A1(_00131_),
    .A2(net3474));
 sg13g2_mux2_1 _08583_ (.A0(_00451_),
    .A1(_00323_),
    .S(net3474),
    .X(_03071_));
 sg13g2_a21oi_1 _08584_ (.A1(net3529),
    .A2(_03071_),
    .Y(_03072_),
    .B1(net3470));
 sg13g2_nor2_1 _08585_ (.A(_00515_),
    .B(net3484),
    .Y(_03073_));
 sg13g2_o21ai_1 _08586_ (.B1(net3521),
    .Y(_03074_),
    .A1(_00419_),
    .A2(net3512));
 sg13g2_mux2_1 _08587_ (.A0(_00163_),
    .A1(_00291_),
    .S(net3485),
    .X(_03075_));
 sg13g2_a21oi_1 _08588_ (.A1(net3537),
    .A2(_03075_),
    .Y(_03076_),
    .B1(net3464));
 sg13g2_o21ai_1 _08589_ (.B1(_03076_),
    .Y(_03077_),
    .A1(_03073_),
    .A2(_03074_));
 sg13g2_a21oi_1 _08590_ (.A1(_03070_),
    .A2(_03072_),
    .Y(_03078_),
    .B1(net3461));
 sg13g2_mux4_1 _08591_ (.S0(net3474),
    .A0(_00227_),
    .A1(_00097_),
    .A2(_00387_),
    .A3(_00259_),
    .S1(net3535),
    .X(_03079_));
 sg13g2_o21ai_1 _08592_ (.B1(net3529),
    .Y(_03080_),
    .A1(net3647),
    .A2(_00355_));
 sg13g2_a21oi_1 _08593_ (.A1(_01715_),
    .A2(net3511),
    .Y(_03081_),
    .B1(_03080_));
 sg13g2_a21oi_1 _08594_ (.A1(_00483_),
    .A2(net3520),
    .Y(_03082_),
    .B1(_03081_));
 sg13g2_o21ai_1 _08595_ (.B1(_02483_),
    .Y(_03083_),
    .A1(_02463_),
    .A2(_03082_));
 sg13g2_a221oi_1 _08596_ (.B2(net3430),
    .C1(_03083_),
    .B1(_03079_),
    .A1(_03077_),
    .Y(_03084_),
    .A2(_03078_));
 sg13g2_nand2b_1 _08597_ (.Y(_03085_),
    .B(net3516),
    .A_N(_00155_));
 sg13g2_a21oi_1 _08598_ (.A1(_01677_),
    .A2(net3479),
    .Y(_03086_),
    .B1(net3531));
 sg13g2_mux2_1 _08599_ (.A0(_00475_),
    .A1(_00347_),
    .S(net3479),
    .X(_03087_));
 sg13g2_a221oi_1 _08600_ (.B2(net3534),
    .C1(net3472),
    .B1(_03087_),
    .A1(_03085_),
    .Y(_03088_),
    .A2(_03086_));
 sg13g2_mux2_1 _08601_ (.A0(_00539_),
    .A1(_00443_),
    .S(net3479),
    .X(_03089_));
 sg13g2_nand2b_1 _08602_ (.Y(_03090_),
    .B(net3646),
    .A_N(_00187_));
 sg13g2_a21oi_1 _08603_ (.A1(_01678_),
    .A2(net3479),
    .Y(_03091_),
    .B1(net3519));
 sg13g2_a221oi_1 _08604_ (.B2(_03091_),
    .C1(net3467),
    .B1(_03090_),
    .A1(net3519),
    .Y(_03092_),
    .A2(_03089_));
 sg13g2_or3_1 _08605_ (.A(net3462),
    .B(_03088_),
    .C(_03092_),
    .X(_03093_));
 sg13g2_mux4_1 _08606_ (.S0(net3478),
    .A0(_00251_),
    .A1(_00121_),
    .A2(_00411_),
    .A3(_00283_),
    .S1(net3531),
    .X(_03094_));
 sg13g2_nand2_1 _08607_ (.Y(_03095_),
    .A(net3431),
    .B(_03094_));
 sg13g2_nand2_1 _08608_ (.Y(_03096_),
    .A(_00507_),
    .B(net3519));
 sg13g2_nor2_1 _08609_ (.A(_00089_),
    .B(net3479),
    .Y(_03097_));
 sg13g2_o21ai_1 _08610_ (.B1(net3534),
    .Y(_03098_),
    .A1(_00379_),
    .A2(net3646));
 sg13g2_o21ai_1 _08611_ (.B1(_03096_),
    .Y(_03099_),
    .A1(_03097_),
    .A2(_03098_));
 sg13g2_a21oi_1 _08612_ (.A1(net3426),
    .A2(_03099_),
    .Y(_03100_),
    .B1(net3386));
 sg13g2_and3_2 _08613_ (.X(_03101_),
    .A(_03093_),
    .B(_03095_),
    .C(_03100_));
 sg13g2_nand2b_1 _08614_ (.Y(_03102_),
    .B(net3515),
    .A_N(_00147_));
 sg13g2_a21oi_1 _08615_ (.A1(_01628_),
    .A2(net3508),
    .Y(_03103_),
    .B1(net3552));
 sg13g2_mux2_1 _08616_ (.A0(_00467_),
    .A1(_00339_),
    .S(net3508),
    .X(_03104_));
 sg13g2_a221oi_1 _08617_ (.B2(net3552),
    .C1(net3472),
    .B1(_03104_),
    .A1(_03102_),
    .Y(_03105_),
    .A2(_03103_));
 sg13g2_nor2_1 _08618_ (.A(_00531_),
    .B(net3508),
    .Y(_03106_));
 sg13g2_a21oi_1 _08619_ (.A1(_01631_),
    .A2(net3508),
    .Y(_03107_),
    .B1(_03106_));
 sg13g2_nand2_1 _08620_ (.Y(_03108_),
    .A(_01632_),
    .B(net3651));
 sg13g2_a21oi_1 _08621_ (.A1(_01633_),
    .A2(net3508),
    .Y(_03109_),
    .B1(net3527));
 sg13g2_a221oi_1 _08622_ (.B2(_03109_),
    .C1(net3468),
    .B1(_03108_),
    .A1(net3526),
    .Y(_03110_),
    .A2(_03107_));
 sg13g2_nand2b_1 _08623_ (.Y(_03111_),
    .B(_02452_),
    .A_N(_03105_));
 sg13g2_mux4_1 _08624_ (.S0(net3507),
    .A0(_00243_),
    .A1(_00113_),
    .A2(_00403_),
    .A3(_00275_),
    .S1(net3551),
    .X(_03112_));
 sg13g2_nand2_1 _08625_ (.Y(_03113_),
    .A(_00499_),
    .B(net3526));
 sg13g2_nor2_1 _08626_ (.A(_00081_),
    .B(net3507),
    .Y(_03114_));
 sg13g2_o21ai_1 _08627_ (.B1(net3551),
    .Y(_03115_),
    .A1(_00371_),
    .A2(net3651));
 sg13g2_o21ai_1 _08628_ (.B1(_03113_),
    .Y(_03116_),
    .A1(_03114_),
    .A2(_03115_));
 sg13g2_a221oi_1 _08629_ (.B2(net3429),
    .C1(net3386),
    .B1(_03116_),
    .A1(net3433),
    .Y(_03117_),
    .A2(_03112_));
 sg13g2_o21ai_1 _08630_ (.B1(_03117_),
    .Y(_03118_),
    .A1(_03110_),
    .A2(_03111_));
 sg13g2_nor2_1 _08631_ (.A(net3234),
    .B(_03118_),
    .Y(_03119_));
 sg13g2_a21oi_2 _08632_ (.B1(_03119_),
    .Y(_03120_),
    .A2(_03101_),
    .A1(net3231));
 sg13g2_nor2_1 _08633_ (.A(net3130),
    .B(_03120_),
    .Y(_03121_));
 sg13g2_a21oi_2 _08634_ (.B1(_03121_),
    .Y(_03122_),
    .A2(_03084_),
    .A1(net3132));
 sg13g2_nor2b_1 _08635_ (.A(_03122_),
    .B_N(net3728),
    .Y(_03123_));
 sg13g2_nand2b_1 _08636_ (.Y(_03124_),
    .B(net3513),
    .A_N(_00139_));
 sg13g2_a21oi_1 _08637_ (.A1(_01587_),
    .A2(net3494),
    .Y(_03125_),
    .B1(net3542));
 sg13g2_nor2_1 _08638_ (.A(_00331_),
    .B(net3512),
    .Y(_03126_));
 sg13g2_a21oi_1 _08639_ (.A1(_01588_),
    .A2(net3513),
    .Y(_03127_),
    .B1(_03126_));
 sg13g2_a221oi_1 _08640_ (.B2(net3542),
    .C1(net3470),
    .B1(_03127_),
    .A1(_03124_),
    .Y(_03128_),
    .A2(_03125_));
 sg13g2_a21oi_1 _08641_ (.A1(_01590_),
    .A2(net3494),
    .Y(_03129_),
    .B1(net3544));
 sg13g2_o21ai_1 _08642_ (.B1(_03129_),
    .Y(_03130_),
    .A1(_00523_),
    .A2(net3494));
 sg13g2_mux2_1 _08643_ (.A0(_00171_),
    .A1(_00299_),
    .S(net3496),
    .X(_03131_));
 sg13g2_a21oi_1 _08644_ (.A1(net3543),
    .A2(_03131_),
    .Y(_03132_),
    .B1(net3464));
 sg13g2_a21o_1 _08645_ (.A2(_03132_),
    .A1(_03130_),
    .B1(net3460),
    .X(_03133_));
 sg13g2_mux4_1 _08646_ (.S0(net3495),
    .A0(_00235_),
    .A1(_00105_),
    .A2(_00395_),
    .A3(_00267_),
    .S1(net3542),
    .X(_03134_));
 sg13g2_nand2_1 _08647_ (.Y(_03135_),
    .A(_00491_),
    .B(net3523));
 sg13g2_nor2_1 _08648_ (.A(_00073_),
    .B(net3495),
    .Y(_03136_));
 sg13g2_o21ai_1 _08649_ (.B1(net3543),
    .Y(_03137_),
    .A1(_00363_),
    .A2(net3648));
 sg13g2_o21ai_1 _08650_ (.B1(_03135_),
    .Y(_03138_),
    .A1(_03136_),
    .A2(_03137_));
 sg13g2_a221oi_1 _08651_ (.B2(net3428),
    .C1(net3386),
    .B1(_03138_),
    .A1(net3432),
    .Y(_03139_),
    .A2(_03134_));
 sg13g2_o21ai_1 _08652_ (.B1(_03139_),
    .Y(_03140_),
    .A1(_03128_),
    .A2(_03133_));
 sg13g2_nor2_1 _08653_ (.A(net3135),
    .B(_03140_),
    .Y(_03141_));
 sg13g2_a21oi_2 _08654_ (.B1(_03141_),
    .Y(_03142_),
    .A2(net3326),
    .A1(net3135));
 sg13g2_a21oi_1 _08655_ (.A1(net3723),
    .A2(net3326),
    .Y(_03143_),
    .B1(net3416));
 sg13g2_o21ai_1 _08656_ (.B1(_03143_),
    .Y(_03144_),
    .A1(net3456),
    .A2(_03120_));
 sg13g2_nor3_1 _08657_ (.A(_03068_),
    .B(_03123_),
    .C(_03144_),
    .Y(_03145_));
 sg13g2_o21ai_1 _08658_ (.B1(_03145_),
    .Y(_03146_),
    .A1(net3725),
    .A2(_03142_));
 sg13g2_mux2_2 _08659_ (.A0(\cpu.PCreg0[4] ),
    .A1(\cpu.PCreg1[4] ),
    .S(net3637),
    .X(\cpu.PC[4] ));
 sg13g2_xnor2_1 _08660_ (.Y(_03147_),
    .A(_01976_),
    .B(_01977_));
 sg13g2_nor2_1 _08661_ (.A(net3406),
    .B(_03147_),
    .Y(_03148_));
 sg13g2_a21oi_2 _08662_ (.B1(_03148_),
    .Y(_03149_),
    .A2(\cpu.PC[4] ),
    .A1(net3406));
 sg13g2_a21o_1 _08663_ (.A2(\cpu.PC[4] ),
    .A1(net3406),
    .B1(_03148_),
    .X(_03150_));
 sg13g2_o21ai_1 _08664_ (.B1(_03146_),
    .Y(_03151_),
    .A1(_02714_),
    .A2(net3124));
 sg13g2_nand2_1 _08665_ (.Y(_03152_),
    .A(\bsq[17] ),
    .B(net3931));
 sg13g2_o21ai_1 _08666_ (.B1(_03152_),
    .Y(uio_out[2]),
    .A1(net3931),
    .A2(_03151_));
 sg13g2_a21oi_1 _08667_ (.A1(net3899),
    .A2(_03151_),
    .Y(_03153_),
    .B1(_02589_));
 sg13g2_o21ai_1 _08668_ (.B1(_03153_),
    .Y(_03154_),
    .A1(net3899),
    .A2(uio_out[2]));
 sg13g2_a21oi_1 _08669_ (.A1(\jtag0.bssh[18] ),
    .A2(net3928),
    .Y(_03155_),
    .B1(net3894));
 sg13g2_a22oi_1 _08670_ (.Y(_01303_),
    .B1(_03154_),
    .B2(_03155_),
    .A2(net3894),
    .A1(_01551_));
 sg13g2_xnor2_1 _08671_ (.Y(_03156_),
    .A(_01840_),
    .B(_02059_));
 sg13g2_mux2_2 _08672_ (.A0(\cpu.PCreg0[11] ),
    .A1(\cpu.PCreg1[11] ),
    .S(net3630),
    .X(\cpu.PC[11] ));
 sg13g2_o21ai_1 _08673_ (.B1(_02622_),
    .Y(_03157_),
    .A1(net3403),
    .A2(\cpu.PC[11] ));
 sg13g2_a21oi_1 _08674_ (.A1(net3402),
    .A2(_03156_),
    .Y(_03158_),
    .B1(_03157_));
 sg13g2_a21oi_1 _08675_ (.A1(_01710_),
    .A2(net3496),
    .Y(_03159_),
    .B1(net3543));
 sg13g2_o21ai_1 _08676_ (.B1(_03159_),
    .Y(_03160_),
    .A1(_00132_),
    .A2(net3496));
 sg13g2_mux2_1 _08677_ (.A0(_00452_),
    .A1(_00324_),
    .S(net3496),
    .X(_03161_));
 sg13g2_a21oi_1 _08678_ (.A1(net3543),
    .A2(_03161_),
    .Y(_03162_),
    .B1(net3473));
 sg13g2_a21oi_1 _08679_ (.A1(_01713_),
    .A2(net3496),
    .Y(_03163_),
    .B1(net3543));
 sg13g2_o21ai_1 _08680_ (.B1(_03163_),
    .Y(_03164_),
    .A1(_00516_),
    .A2(net3496));
 sg13g2_mux2_1 _08681_ (.A0(_00164_),
    .A1(_00292_),
    .S(net3496),
    .X(_03165_));
 sg13g2_a21oi_1 _08682_ (.A1(net3543),
    .A2(_03165_),
    .Y(_03166_),
    .B1(net3464));
 sg13g2_nand2_1 _08683_ (.Y(_03167_),
    .A(_03164_),
    .B(_03166_));
 sg13g2_a21oi_1 _08684_ (.A1(_03160_),
    .A2(_03162_),
    .Y(_03168_),
    .B1(net3460));
 sg13g2_mux4_1 _08685_ (.S0(net3493),
    .A0(_00228_),
    .A1(_00098_),
    .A2(_00388_),
    .A3(_00260_),
    .S1(net3541),
    .X(_03169_));
 sg13g2_and2_1 _08686_ (.A(_00484_),
    .B(net3523),
    .X(_03170_));
 sg13g2_mux2_1 _08687_ (.A0(_00066_),
    .A1(_00356_),
    .S(net3496),
    .X(_03171_));
 sg13g2_a21oi_1 _08688_ (.A1(net3543),
    .A2(_03171_),
    .Y(_03172_),
    .B1(_03170_));
 sg13g2_o21ai_1 _08689_ (.B1(_02483_),
    .Y(_03173_),
    .A1(_02463_),
    .A2(_03172_));
 sg13g2_a221oi_1 _08690_ (.B2(net3432),
    .C1(_03173_),
    .B1(_03169_),
    .A1(_03167_),
    .Y(_03174_),
    .A2(_03168_));
 sg13g2_nand2b_1 _08691_ (.Y(_03175_),
    .B(net3515),
    .A_N(_00148_));
 sg13g2_a21oi_1 _08692_ (.A1(_01634_),
    .A2(net3503),
    .Y(_03176_),
    .B1(net3547));
 sg13g2_mux2_1 _08693_ (.A0(_00468_),
    .A1(_00340_),
    .S(net3503),
    .X(_03177_));
 sg13g2_a221oi_1 _08694_ (.B2(net3547),
    .C1(net3472),
    .B1(_03177_),
    .A1(_03175_),
    .Y(_03178_),
    .A2(_03176_));
 sg13g2_mux2_1 _08695_ (.A0(_00532_),
    .A1(_00436_),
    .S(net3501),
    .X(_03179_));
 sg13g2_nand2_1 _08696_ (.Y(_03180_),
    .A(_01637_),
    .B(net3651));
 sg13g2_a21oi_1 _08697_ (.A1(_01638_),
    .A2(net3501),
    .Y(_03181_),
    .B1(net3525));
 sg13g2_a221oi_1 _08698_ (.B2(_03181_),
    .C1(net3466),
    .B1(_03180_),
    .A1(net3525),
    .Y(_03182_),
    .A2(_03179_));
 sg13g2_or3_1 _08699_ (.A(net3463),
    .B(_03178_),
    .C(_03182_),
    .X(_03183_));
 sg13g2_mux4_1 _08700_ (.S0(net3500),
    .A0(_00244_),
    .A1(_00114_),
    .A2(_00404_),
    .A3(_00276_),
    .S1(net3546),
    .X(_03184_));
 sg13g2_nand2_1 _08701_ (.Y(_03185_),
    .A(net3433),
    .B(_03184_));
 sg13g2_nand2_1 _08702_ (.Y(_03186_),
    .A(_00500_),
    .B(net3524));
 sg13g2_nor2_1 _08703_ (.A(_00082_),
    .B(net3500),
    .Y(_03187_));
 sg13g2_o21ai_1 _08704_ (.B1(net3546),
    .Y(_03188_),
    .A1(_00372_),
    .A2(net3649));
 sg13g2_o21ai_1 _08705_ (.B1(_03186_),
    .Y(_03189_),
    .A1(_03187_),
    .A2(_03188_));
 sg13g2_a21oi_1 _08706_ (.A1(net3427),
    .A2(_03189_),
    .Y(_03190_),
    .B1(net3386));
 sg13g2_nand3_1 _08707_ (.B(_03185_),
    .C(_03190_),
    .A(_03183_),
    .Y(_03191_));
 sg13g2_nor2_1 _08708_ (.A(net3234),
    .B(_03191_),
    .Y(_03192_));
 sg13g2_a21oi_2 _08709_ (.B1(_03192_),
    .Y(_03193_),
    .A2(net3234),
    .A1(_02469_));
 sg13g2_nor2_1 _08710_ (.A(net3132),
    .B(_03193_),
    .Y(_03194_));
 sg13g2_a21oi_2 _08711_ (.B1(_03194_),
    .Y(_03195_),
    .A2(_03174_),
    .A1(net3132));
 sg13g2_nor2b_1 _08712_ (.A(_03195_),
    .B_N(net3728),
    .Y(_03196_));
 sg13g2_nand2b_1 _08713_ (.Y(_03197_),
    .B(net3514),
    .A_N(_00140_));
 sg13g2_a21oi_1 _08714_ (.A1(_01591_),
    .A2(net3506),
    .Y(_03198_),
    .B1(net3550));
 sg13g2_nor2_1 _08715_ (.A(_00332_),
    .B(net3514),
    .Y(_03199_));
 sg13g2_a21oi_1 _08716_ (.A1(_01592_),
    .A2(net3514),
    .Y(_03200_),
    .B1(_03199_));
 sg13g2_a221oi_1 _08717_ (.B2(net3550),
    .C1(net3471),
    .B1(_03200_),
    .A1(_03197_),
    .Y(_03201_),
    .A2(_03198_));
 sg13g2_nor2_1 _08718_ (.A(_00524_),
    .B(net3505),
    .Y(_03202_));
 sg13g2_o21ai_1 _08719_ (.B1(net3527),
    .Y(_03203_),
    .A1(_00428_),
    .A2(net3514));
 sg13g2_o21ai_1 _08720_ (.B1(net3550),
    .Y(_03204_),
    .A1(_00300_),
    .A2(net3514));
 sg13g2_a21oi_1 _08721_ (.A1(_01595_),
    .A2(net3650),
    .Y(_03205_),
    .B1(_03204_));
 sg13g2_o21ai_1 _08722_ (.B1(net3471),
    .Y(_03206_),
    .A1(_03202_),
    .A2(_03203_));
 sg13g2_o21ai_1 _08723_ (.B1(_02452_),
    .Y(_03207_),
    .A1(_03205_),
    .A2(_03206_));
 sg13g2_mux4_1 _08724_ (.S0(net3506),
    .A0(_00236_),
    .A1(_00106_),
    .A2(_00396_),
    .A3(_00268_),
    .S1(net3550),
    .X(_03208_));
 sg13g2_nand2_1 _08725_ (.Y(_03209_),
    .A(_00492_),
    .B(net3527));
 sg13g2_nor2_1 _08726_ (.A(_00074_),
    .B(net3506),
    .Y(_03210_));
 sg13g2_o21ai_1 _08727_ (.B1(net3550),
    .Y(_03211_),
    .A1(_00364_),
    .A2(net3650));
 sg13g2_o21ai_1 _08728_ (.B1(_03209_),
    .Y(_03212_),
    .A1(_03210_),
    .A2(_03211_));
 sg13g2_a221oi_1 _08729_ (.B2(net3429),
    .C1(_02482_),
    .B1(_03212_),
    .A1(net3433),
    .Y(_03213_),
    .A2(_03208_));
 sg13g2_o21ai_1 _08730_ (.B1(_03213_),
    .Y(_03214_),
    .A1(_03201_),
    .A2(_03207_));
 sg13g2_nor2_1 _08731_ (.A(net3136),
    .B(_03214_),
    .Y(_03215_));
 sg13g2_a21oi_2 _08732_ (.B1(_03215_),
    .Y(_03216_),
    .A2(net3136),
    .A1(_02469_));
 sg13g2_a21oi_1 _08733_ (.A1(_02469_),
    .A2(net3723),
    .Y(_03217_),
    .B1(net3416));
 sg13g2_o21ai_1 _08734_ (.B1(_03217_),
    .Y(_03218_),
    .A1(net3456),
    .A2(_03193_));
 sg13g2_nor3_1 _08735_ (.A(_03158_),
    .B(_03196_),
    .C(_03218_),
    .Y(_03219_));
 sg13g2_o21ai_1 _08736_ (.B1(_03219_),
    .Y(_03220_),
    .A1(net3725),
    .A2(_03216_));
 sg13g2_mux2_2 _08737_ (.A0(\cpu.PCreg0[3] ),
    .A1(\cpu.PCreg1[3] ),
    .S(net3636),
    .X(\cpu.PC[3] ));
 sg13g2_nor2_1 _08738_ (.A(net3405),
    .B(\cpu.PC[3] ),
    .Y(_03221_));
 sg13g2_xnor2_1 _08739_ (.Y(_03222_),
    .A(_01974_),
    .B(_01975_));
 sg13g2_a21oi_2 _08740_ (.B1(_03221_),
    .Y(_03223_),
    .A2(_03222_),
    .A1(net3405));
 sg13g2_inv_1 _08741_ (.Y(_03224_),
    .A(_03223_));
 sg13g2_o21ai_1 _08742_ (.B1(_03220_),
    .Y(_03225_),
    .A1(_02714_),
    .A2(_03223_));
 sg13g2_nand2_1 _08743_ (.Y(_03226_),
    .A(\bsq[16] ),
    .B(net3931));
 sg13g2_o21ai_1 _08744_ (.B1(_03226_),
    .Y(uio_out[1]),
    .A1(net3929),
    .A2(_03225_));
 sg13g2_a21oi_1 _08745_ (.A1(net3899),
    .A2(_03225_),
    .Y(_03227_),
    .B1(_02589_));
 sg13g2_o21ai_1 _08746_ (.B1(_03227_),
    .Y(_03228_),
    .A1(net3899),
    .A2(uio_out[1]));
 sg13g2_a21oi_1 _08747_ (.A1(\jtag0.bssh[17] ),
    .A2(net3928),
    .Y(_03229_),
    .B1(net3894));
 sg13g2_a22oi_1 _08748_ (.Y(_01302_),
    .B1(_03228_),
    .B2(_03229_),
    .A2(net3894),
    .A1(_01552_));
 sg13g2_xnor2_1 _08749_ (.Y(_03230_),
    .A(_02038_),
    .B(_02056_));
 sg13g2_mux2_2 _08750_ (.A0(\cpu.PCreg0[10] ),
    .A1(\cpu.PCreg1[10] ),
    .S(net3635),
    .X(\cpu.PC[10] ));
 sg13g2_o21ai_1 _08751_ (.B1(_02622_),
    .Y(_03231_),
    .A1(net3402),
    .A2(\cpu.PC[10] ));
 sg13g2_a21oi_1 _08752_ (.A1(net3403),
    .A2(_03230_),
    .Y(_03232_),
    .B1(_03231_));
 sg13g2_a21oi_1 _08753_ (.A1(_01708_),
    .A2(net3485),
    .Y(_03233_),
    .B1(net3537));
 sg13g2_o21ai_1 _08754_ (.B1(_03233_),
    .Y(_03234_),
    .A1(_00133_),
    .A2(net3485));
 sg13g2_mux2_1 _08755_ (.A0(_00453_),
    .A1(_00325_),
    .S(net3485),
    .X(_03235_));
 sg13g2_a21oi_1 _08756_ (.A1(net3537),
    .A2(_03235_),
    .Y(_03236_),
    .B1(net3469));
 sg13g2_nor2_1 _08757_ (.A(_00517_),
    .B(net3486),
    .Y(_03237_));
 sg13g2_o21ai_1 _08758_ (.B1(net3521),
    .Y(_03238_),
    .A1(_00421_),
    .A2(net3512));
 sg13g2_mux2_1 _08759_ (.A0(_00165_),
    .A1(_00293_),
    .S(net3486),
    .X(_03239_));
 sg13g2_a21oi_1 _08760_ (.A1(net3536),
    .A2(_03239_),
    .Y(_03240_),
    .B1(net3464));
 sg13g2_o21ai_1 _08761_ (.B1(_03240_),
    .Y(_03241_),
    .A1(_03237_),
    .A2(_03238_));
 sg13g2_a21oi_1 _08762_ (.A1(_03234_),
    .A2(_03236_),
    .Y(_03242_),
    .B1(net3460));
 sg13g2_mux4_1 _08763_ (.S0(net3486),
    .A0(_00229_),
    .A1(_00099_),
    .A2(_00389_),
    .A3(_00261_),
    .S1(net3536),
    .X(_03243_));
 sg13g2_and2_1 _08764_ (.A(_00485_),
    .B(net3523),
    .X(_03244_));
 sg13g2_mux2_1 _08765_ (.A0(_00067_),
    .A1(_00357_),
    .S(net3487),
    .X(_03245_));
 sg13g2_a21oi_1 _08766_ (.A1(net3539),
    .A2(_03245_),
    .Y(_03246_),
    .B1(_03244_));
 sg13g2_o21ai_1 _08767_ (.B1(_02483_),
    .Y(_03247_),
    .A1(_02463_),
    .A2(_03246_));
 sg13g2_a221oi_1 _08768_ (.B2(net3432),
    .C1(_03247_),
    .B1(_03243_),
    .A1(_03241_),
    .Y(_03248_),
    .A2(_03242_));
 sg13g2_nand2b_1 _08769_ (.Y(_03249_),
    .B(net3514),
    .A_N(_00149_));
 sg13g2_a21oi_1 _08770_ (.A1(_01639_),
    .A2(net3509),
    .Y(_03250_),
    .B1(net3551));
 sg13g2_mux2_1 _08771_ (.A0(_00469_),
    .A1(_00341_),
    .S(net3508),
    .X(_03251_));
 sg13g2_a221oi_1 _08772_ (.B2(net3551),
    .C1(net3471),
    .B1(_03251_),
    .A1(_03249_),
    .Y(_03252_),
    .A2(_03250_));
 sg13g2_nor2_1 _08773_ (.A(_00533_),
    .B(net3508),
    .Y(_03253_));
 sg13g2_a21oi_1 _08774_ (.A1(_01642_),
    .A2(net3508),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_nand2_1 _08775_ (.Y(_03255_),
    .A(_01643_),
    .B(net3650));
 sg13g2_a21oi_1 _08776_ (.A1(_01644_),
    .A2(net3507),
    .Y(_03256_),
    .B1(net3526));
 sg13g2_a221oi_1 _08777_ (.B2(_03256_),
    .C1(net3466),
    .B1(_03255_),
    .A1(net3526),
    .Y(_03257_),
    .A2(_03254_));
 sg13g2_nand2b_1 _08778_ (.Y(_03258_),
    .B(_02452_),
    .A_N(_03252_));
 sg13g2_mux4_1 _08779_ (.S0(net3501),
    .A0(_00245_),
    .A1(_00115_),
    .A2(_00405_),
    .A3(_00277_),
    .S1(net3548),
    .X(_03259_));
 sg13g2_nand2_1 _08780_ (.Y(_03260_),
    .A(_00501_),
    .B(net3525));
 sg13g2_nor2_1 _08781_ (.A(_00083_),
    .B(net3502),
    .Y(_03261_));
 sg13g2_o21ai_1 _08782_ (.B1(net3548),
    .Y(_03262_),
    .A1(_00373_),
    .A2(net3649));
 sg13g2_o21ai_1 _08783_ (.B1(_03260_),
    .Y(_03263_),
    .A1(_03261_),
    .A2(_03262_));
 sg13g2_a221oi_1 _08784_ (.B2(net3427),
    .C1(_02482_),
    .B1(_03263_),
    .A1(net3433),
    .Y(_03264_),
    .A2(_03259_));
 sg13g2_o21ai_1 _08785_ (.B1(_03264_),
    .Y(_03265_),
    .A1(_03257_),
    .A2(_03258_));
 sg13g2_nor2_1 _08786_ (.A(net3233),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_a21oi_2 _08787_ (.B1(_03266_),
    .Y(_03267_),
    .A2(net3233),
    .A1(_02498_));
 sg13g2_nor2_1 _08788_ (.A(net3133),
    .B(_03267_),
    .Y(_03268_));
 sg13g2_a21oi_2 _08789_ (.B1(_03268_),
    .Y(_03269_),
    .A2(_03248_),
    .A1(net3133));
 sg13g2_nor2b_1 _08790_ (.A(_03269_),
    .B_N(net3728),
    .Y(_03270_));
 sg13g2_mux2_1 _08791_ (.A0(_00141_),
    .A1(_00205_),
    .S(net3482),
    .X(_03271_));
 sg13g2_nand2b_1 _08792_ (.Y(_03272_),
    .B(net3482),
    .A_N(_00333_));
 sg13g2_a21oi_1 _08793_ (.A1(_01596_),
    .A2(net3653),
    .Y(_03273_),
    .B1(net3518));
 sg13g2_a221oi_1 _08794_ (.B2(_03273_),
    .C1(net3472),
    .B1(_03272_),
    .A1(net3518),
    .Y(_03274_),
    .A2(_03271_));
 sg13g2_mux2_1 _08795_ (.A0(_00525_),
    .A1(_00429_),
    .S(net3482),
    .X(_03275_));
 sg13g2_nand2_1 _08796_ (.Y(_03276_),
    .A(_01597_),
    .B(net3653));
 sg13g2_a21oi_1 _08797_ (.A1(_01598_),
    .A2(net3482),
    .Y(_03277_),
    .B1(net3518));
 sg13g2_a221oi_1 _08798_ (.B2(_03277_),
    .C1(net3467),
    .B1(_03276_),
    .A1(net3518),
    .Y(_03278_),
    .A2(_03275_));
 sg13g2_or3_1 _08799_ (.A(net3462),
    .B(_03274_),
    .C(_03278_),
    .X(_03279_));
 sg13g2_mux4_1 _08800_ (.S0(net3482),
    .A0(_00237_),
    .A1(_00107_),
    .A2(_00397_),
    .A3(_00269_),
    .S1(net3533),
    .X(_03280_));
 sg13g2_nand2_1 _08801_ (.Y(_03281_),
    .A(net3431),
    .B(_03280_));
 sg13g2_nand2_1 _08802_ (.Y(_03282_),
    .A(_00493_),
    .B(net3520));
 sg13g2_nor2_1 _08803_ (.A(_00075_),
    .B(net3482),
    .Y(_03283_));
 sg13g2_o21ai_1 _08804_ (.B1(net3532),
    .Y(_03284_),
    .A1(_00365_),
    .A2(net3646));
 sg13g2_o21ai_1 _08805_ (.B1(_03282_),
    .Y(_03285_),
    .A1(_03283_),
    .A2(_03284_));
 sg13g2_a21oi_1 _08806_ (.A1(net3426),
    .A2(_03285_),
    .Y(_03286_),
    .B1(net3386));
 sg13g2_and4_2 _08807_ (.A(_02505_),
    .B(_03279_),
    .C(_03281_),
    .D(_03286_),
    .X(_03287_));
 sg13g2_a21oi_2 _08808_ (.B1(_03287_),
    .Y(_03288_),
    .A2(net3139),
    .A1(_02498_));
 sg13g2_a21oi_1 _08809_ (.A1(_02498_),
    .A2(net3723),
    .Y(_03289_),
    .B1(net3416));
 sg13g2_o21ai_1 _08810_ (.B1(_03289_),
    .Y(_03290_),
    .A1(net3456),
    .A2(_03267_));
 sg13g2_nor3_1 _08811_ (.A(_03232_),
    .B(_03270_),
    .C(_03290_),
    .Y(_03291_));
 sg13g2_o21ai_1 _08812_ (.B1(_03291_),
    .Y(_03292_),
    .A1(net3726),
    .A2(_03288_));
 sg13g2_o21ai_1 _08813_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net3142),
    .A2(_02714_));
 sg13g2_nand2_1 _08814_ (.Y(_03294_),
    .A(\bsq[15] ),
    .B(net3932));
 sg13g2_o21ai_1 _08815_ (.B1(_03294_),
    .Y(uio_out[0]),
    .A1(net3932),
    .A2(_03293_));
 sg13g2_a21oi_1 _08816_ (.A1(net3902),
    .A2(_03293_),
    .Y(_03295_),
    .B1(_02589_));
 sg13g2_o21ai_1 _08817_ (.B1(_03295_),
    .Y(_03296_),
    .A1(net3899),
    .A2(uio_out[0]));
 sg13g2_a21oi_1 _08818_ (.A1(\jtag0.bssh[16] ),
    .A2(net3928),
    .Y(_03297_),
    .B1(net3894));
 sg13g2_a22oi_1 _08819_ (.Y(_01301_),
    .B1(_03296_),
    .B2(_03297_),
    .A2(net3897),
    .A1(_01553_));
 sg13g2_nor2_1 _08820_ (.A(net16),
    .B(net3902),
    .Y(_03298_));
 sg13g2_mux2_2 _08821_ (.A0(net16),
    .A1(\bsq[14] ),
    .S(net3934),
    .X(_03299_));
 sg13g2_o21ai_1 _08822_ (.B1(net3731),
    .Y(_03300_),
    .A1(net3736),
    .A2(_03299_));
 sg13g2_a22oi_1 _08823_ (.Y(_03301_),
    .B1(net3882),
    .B2(\jtag0.bssh[15] ),
    .A2(net3895),
    .A1(\jtag0.bssh[14] ));
 sg13g2_o21ai_1 _08824_ (.B1(_03301_),
    .Y(_01300_),
    .A1(_03298_),
    .A2(_03300_));
 sg13g2_mux2_2 _08825_ (.A0(net15),
    .A1(\bsq[13] ),
    .S(net3932),
    .X(_03302_));
 sg13g2_nor2_1 _08826_ (.A(net15),
    .B(net3902),
    .Y(_03303_));
 sg13g2_o21ai_1 _08827_ (.B1(net3731),
    .Y(_03304_),
    .A1(net3736),
    .A2(_03302_));
 sg13g2_a22oi_1 _08828_ (.Y(_03305_),
    .B1(net3882),
    .B2(\jtag0.bssh[14] ),
    .A2(net3895),
    .A1(\jtag0.bssh[13] ));
 sg13g2_o21ai_1 _08829_ (.B1(_03305_),
    .Y(_01299_),
    .A1(_03303_),
    .A2(_03304_));
 sg13g2_nor2_1 _08830_ (.A(net3932),
    .B(net14),
    .Y(_03306_));
 sg13g2_nand2b_1 _08831_ (.Y(_03307_),
    .B(net3932),
    .A_N(\bsq[12] ));
 sg13g2_nor2b_1 _08832_ (.A(_03306_),
    .B_N(_03307_),
    .Y(_03308_));
 sg13g2_nand2b_2 _08833_ (.Y(_03309_),
    .B(_03307_),
    .A_N(_03306_));
 sg13g2_nand2_1 _08834_ (.Y(_03310_),
    .A(net3902),
    .B(_03309_));
 sg13g2_o21ai_1 _08835_ (.B1(_03310_),
    .Y(_03311_),
    .A1(net14),
    .A2(net3902));
 sg13g2_a22oi_1 _08836_ (.Y(_03312_),
    .B1(net3884),
    .B2(\jtag0.bssh[13] ),
    .A2(net3897),
    .A1(\jtag0.bssh[12] ));
 sg13g2_o21ai_1 _08837_ (.B1(_03312_),
    .Y(_01298_),
    .A1(_02589_),
    .A2(_03311_));
 sg13g2_nor2_1 _08838_ (.A(net13),
    .B(net3901),
    .Y(_03313_));
 sg13g2_mux2_2 _08839_ (.A0(net13),
    .A1(\bsq[11] ),
    .S(net3933),
    .X(_03314_));
 sg13g2_o21ai_1 _08840_ (.B1(net3731),
    .Y(_03315_),
    .A1(net3736),
    .A2(_03314_));
 sg13g2_a22oi_1 _08841_ (.Y(_03316_),
    .B1(net3882),
    .B2(\jtag0.bssh[12] ),
    .A2(net3895),
    .A1(\jtag0.bssh[11] ));
 sg13g2_o21ai_1 _08842_ (.B1(_03316_),
    .Y(_01297_),
    .A1(_03313_),
    .A2(_03315_));
 sg13g2_mux2_2 _08843_ (.A0(net12),
    .A1(\bsq[10] ),
    .S(net3933),
    .X(_03317_));
 sg13g2_nor2_1 _08844_ (.A(net12),
    .B(net3901),
    .Y(_03318_));
 sg13g2_o21ai_1 _08845_ (.B1(net3732),
    .Y(_03319_),
    .A1(net3736),
    .A2(_03317_));
 sg13g2_a22oi_1 _08846_ (.Y(_03320_),
    .B1(net3882),
    .B2(\jtag0.bssh[11] ),
    .A2(net3895),
    .A1(\jtag0.bssh[10] ));
 sg13g2_o21ai_1 _08847_ (.B1(_03320_),
    .Y(_01296_),
    .A1(_03318_),
    .A2(_03319_));
 sg13g2_mux2_2 _08848_ (.A0(net11),
    .A1(\bsq[9] ),
    .S(net3934),
    .X(_03321_));
 sg13g2_nor2_1 _08849_ (.A(net11),
    .B(net3901),
    .Y(_03322_));
 sg13g2_o21ai_1 _08850_ (.B1(net3732),
    .Y(_03323_),
    .A1(net3736),
    .A2(_03321_));
 sg13g2_a22oi_1 _08851_ (.Y(_03324_),
    .B1(net3882),
    .B2(\jtag0.bssh[10] ),
    .A2(net3895),
    .A1(\jtag0.bssh[9] ));
 sg13g2_o21ai_1 _08852_ (.B1(_03324_),
    .Y(_01295_),
    .A1(_03322_),
    .A2(_03323_));
 sg13g2_mux2_2 _08853_ (.A0(net10),
    .A1(\bsq[8] ),
    .S(net3933),
    .X(_03325_));
 sg13g2_nor2_1 _08854_ (.A(net10),
    .B(net3901),
    .Y(_03326_));
 sg13g2_o21ai_1 _08855_ (.B1(net3732),
    .Y(_03327_),
    .A1(net3736),
    .A2(_03325_));
 sg13g2_a22oi_1 _08856_ (.Y(_03328_),
    .B1(net3883),
    .B2(\jtag0.bssh[9] ),
    .A2(net3896),
    .A1(\jtag0.bssh[8] ));
 sg13g2_o21ai_1 _08857_ (.B1(_03328_),
    .Y(_01294_),
    .A1(_03326_),
    .A2(_03327_));
 sg13g2_mux2_2 _08858_ (.A0(net9),
    .A1(\bsq[7] ),
    .S(net3933),
    .X(_03329_));
 sg13g2_nor2_1 _08859_ (.A(net9),
    .B(net3903),
    .Y(_03330_));
 sg13g2_o21ai_1 _08860_ (.B1(net3731),
    .Y(_03331_),
    .A1(net3736),
    .A2(_03329_));
 sg13g2_a22oi_1 _08861_ (.Y(_03332_),
    .B1(net3882),
    .B2(\jtag0.bssh[8] ),
    .A2(net3895),
    .A1(\jtag0.bssh[7] ));
 sg13g2_o21ai_1 _08862_ (.B1(_03332_),
    .Y(_01293_),
    .A1(_03330_),
    .A2(_03331_));
 sg13g2_mux2_2 _08863_ (.A0(net8),
    .A1(\bsq[6] ),
    .S(net3933),
    .X(_03333_));
 sg13g2_nor2_1 _08864_ (.A(net8),
    .B(net3903),
    .Y(_03334_));
 sg13g2_o21ai_1 _08865_ (.B1(net3732),
    .Y(_03335_),
    .A1(net3737),
    .A2(_03333_));
 sg13g2_a22oi_1 _08866_ (.Y(_03336_),
    .B1(net3882),
    .B2(\jtag0.bssh[7] ),
    .A2(net3895),
    .A1(\jtag0.bssh[6] ));
 sg13g2_o21ai_1 _08867_ (.B1(_03336_),
    .Y(_01292_),
    .A1(_03334_),
    .A2(_03335_));
 sg13g2_mux2_2 _08868_ (.A0(net7),
    .A1(\bsq[5] ),
    .S(net3933),
    .X(_03337_));
 sg13g2_nor2_1 _08869_ (.A(net7),
    .B(net3901),
    .Y(_03338_));
 sg13g2_o21ai_1 _08870_ (.B1(net3731),
    .Y(_03339_),
    .A1(net3737),
    .A2(_03337_));
 sg13g2_a22oi_1 _08871_ (.Y(_03340_),
    .B1(net3883),
    .B2(\jtag0.bssh[6] ),
    .A2(net3896),
    .A1(\jtag0.bssh[5] ));
 sg13g2_o21ai_1 _08872_ (.B1(_03340_),
    .Y(_01291_),
    .A1(_03338_),
    .A2(_03339_));
 sg13g2_mux2_2 _08873_ (.A0(net6),
    .A1(\bsq[4] ),
    .S(net3930),
    .X(_03341_));
 sg13g2_nor2_1 _08874_ (.A(net6),
    .B(net3901),
    .Y(_03342_));
 sg13g2_o21ai_1 _08875_ (.B1(net3730),
    .Y(_03343_),
    .A1(net3734),
    .A2(_03341_));
 sg13g2_a22oi_1 _08876_ (.Y(_03344_),
    .B1(net3883),
    .B2(\jtag0.bssh[5] ),
    .A2(net3894),
    .A1(\jtag0.bssh[4] ));
 sg13g2_o21ai_1 _08877_ (.B1(_03344_),
    .Y(_01290_),
    .A1(_03342_),
    .A2(_03343_));
 sg13g2_mux2_1 _08878_ (.A0(net5),
    .A1(\bsq[3] ),
    .S(net3929),
    .X(_03345_));
 sg13g2_nor2_1 _08879_ (.A(net5),
    .B(net3899),
    .Y(_03346_));
 sg13g2_o21ai_1 _08880_ (.B1(net3729),
    .Y(_03347_),
    .A1(net3734),
    .A2(_03345_));
 sg13g2_a22oi_1 _08881_ (.Y(_03348_),
    .B1(net3884),
    .B2(\jtag0.bssh[4] ),
    .A2(net3897),
    .A1(\jtag0.bssh[3] ));
 sg13g2_o21ai_1 _08882_ (.B1(_03348_),
    .Y(_01289_),
    .A1(_03346_),
    .A2(_03347_));
 sg13g2_mux2_1 _08883_ (.A0(net4),
    .A1(\bsq[2] ),
    .S(net3929),
    .X(rxd));
 sg13g2_nor2_1 _08884_ (.A(net4),
    .B(net3899),
    .Y(_03349_));
 sg13g2_o21ai_1 _08885_ (.B1(net3729),
    .Y(_03350_),
    .A1(net3734),
    .A2(rxd));
 sg13g2_a22oi_1 _08886_ (.Y(_03351_),
    .B1(net3884),
    .B2(\jtag0.bssh[3] ),
    .A2(net3897),
    .A1(\jtag0.bssh[2] ));
 sg13g2_o21ai_1 _08887_ (.B1(_03351_),
    .Y(_01288_),
    .A1(_03349_),
    .A2(_03350_));
 sg13g2_nor2_1 _08888_ (.A(clknet_1_0__leaf_clk),
    .B(net3899),
    .Y(_03352_));
 sg13g2_o21ai_1 _08889_ (.B1(net3729),
    .Y(_03353_),
    .A1(net3734),
    .A2(clknet_1_0__leaf_jclk));
 sg13g2_a22oi_1 _08890_ (.Y(_03354_),
    .B1(net3885),
    .B2(\jtag0.bssh[2] ),
    .A2(net3893),
    .A1(\jtag0.bssh[1] ));
 sg13g2_o21ai_1 _08891_ (.B1(_03354_),
    .Y(_01287_),
    .A1(_03352_),
    .A2(_03353_));
 sg13g2_o21ai_1 _08892_ (.B1(net3953),
    .Y(_03355_),
    .A1(\bsq[0] ),
    .A2(_02565_));
 sg13g2_inv_1 _08893_ (.Y(_00027_),
    .A(net3875));
 sg13g2_a21oi_1 _08894_ (.A1(_01573_),
    .A2(net3953),
    .Y(_03356_),
    .B1(_02589_));
 sg13g2_nor2b_1 _08895_ (.A(\jtag0.bssh[1] ),
    .B_N(net3885),
    .Y(_03357_));
 sg13g2_a221oi_1 _08896_ (.B2(_03356_),
    .C1(_03357_),
    .B1(net3876),
    .A1(_01554_),
    .Y(_01286_),
    .A2(net3893));
 sg13g2_a22oi_1 _08897_ (.Y(_03358_),
    .B1(net3886),
    .B2(\jtag0.stdi ),
    .A2(net3891),
    .A1(\jtag0.idr[31] ));
 sg13g2_inv_1 _08898_ (.Y(_01285_),
    .A(_03358_));
 sg13g2_a22oi_1 _08899_ (.Y(_03359_),
    .B1(net3881),
    .B2(\jtag0.idr[31] ),
    .A2(net3891),
    .A1(\jtag0.idr[30] ));
 sg13g2_inv_1 _08900_ (.Y(_01284_),
    .A(_03359_));
 sg13g2_a22oi_1 _08901_ (.Y(_03360_),
    .B1(net3881),
    .B2(\jtag0.idr[30] ),
    .A2(net3891),
    .A1(\jtag0.idr[29] ));
 sg13g2_inv_1 _08902_ (.Y(_01283_),
    .A(_03360_));
 sg13g2_a22oi_1 _08903_ (.Y(_03361_),
    .B1(net3881),
    .B2(\jtag0.idr[29] ),
    .A2(net3891),
    .A1(\jtag0.idr[28] ));
 sg13g2_inv_1 _08904_ (.Y(_01282_),
    .A(_03361_));
 sg13g2_a22oi_1 _08905_ (.Y(_03362_),
    .B1(net3879),
    .B2(\jtag0.idr[28] ),
    .A2(net3889),
    .A1(\jtag0.idr[27] ));
 sg13g2_inv_1 _08906_ (.Y(_01281_),
    .A(_03362_));
 sg13g2_a22oi_1 _08907_ (.Y(_03363_),
    .B1(net3879),
    .B2(\jtag0.idr[27] ),
    .A2(net3889),
    .A1(\jtag0.idr[26] ));
 sg13g2_inv_1 _08908_ (.Y(_01280_),
    .A(_03363_));
 sg13g2_a22oi_1 _08909_ (.Y(_03364_),
    .B1(net3879),
    .B2(\jtag0.idr[26] ),
    .A2(net3889),
    .A1(\jtag0.idr[25] ));
 sg13g2_inv_1 _08910_ (.Y(_01279_),
    .A(_03364_));
 sg13g2_a22oi_1 _08911_ (.Y(_03365_),
    .B1(net3881),
    .B2(\jtag0.idr[25] ),
    .A2(net3890),
    .A1(\jtag0.idr[24] ));
 sg13g2_inv_1 _08912_ (.Y(_01278_),
    .A(_03365_));
 sg13g2_a22oi_1 _08913_ (.Y(_03366_),
    .B1(net3881),
    .B2(\jtag0.idr[24] ),
    .A2(net3898),
    .A1(\jtag0.idr[23] ));
 sg13g2_inv_1 _08914_ (.Y(_01277_),
    .A(_03366_));
 sg13g2_a22oi_1 _08915_ (.Y(_03367_),
    .B1(net3880),
    .B2(\jtag0.idr[23] ),
    .A2(net3890),
    .A1(\jtag0.idr[22] ));
 sg13g2_inv_1 _08916_ (.Y(_01276_),
    .A(_03367_));
 sg13g2_a22oi_1 _08917_ (.Y(_03368_),
    .B1(net3879),
    .B2(\jtag0.idr[22] ),
    .A2(net3889),
    .A1(\jtag0.idr[21] ));
 sg13g2_inv_1 _08918_ (.Y(_01275_),
    .A(_03368_));
 sg13g2_a22oi_1 _08919_ (.Y(_03369_),
    .B1(net3879),
    .B2(\jtag0.idr[21] ),
    .A2(net3889),
    .A1(\jtag0.idr[20] ));
 sg13g2_inv_1 _08920_ (.Y(_01274_),
    .A(_03369_));
 sg13g2_a22oi_1 _08921_ (.Y(_03370_),
    .B1(net3879),
    .B2(\jtag0.idr[20] ),
    .A2(net3889),
    .A1(\jtag0.idr[19] ));
 sg13g2_inv_1 _08922_ (.Y(_01273_),
    .A(_03370_));
 sg13g2_a22oi_1 _08923_ (.Y(_01272_),
    .B1(net3877),
    .B2(_01555_),
    .A2(net3887),
    .A1(_01556_));
 sg13g2_a22oi_1 _08924_ (.Y(_03371_),
    .B1(net3877),
    .B2(\jtag0.idr[18] ),
    .A2(net3887),
    .A1(\jtag0.idr[17] ));
 sg13g2_inv_1 _08925_ (.Y(_01271_),
    .A(_03371_));
 sg13g2_a22oi_1 _08926_ (.Y(_03372_),
    .B1(net3877),
    .B2(\jtag0.idr[17] ),
    .A2(net3887),
    .A1(\jtag0.idr[16] ));
 sg13g2_inv_1 _08927_ (.Y(_01270_),
    .A(_03372_));
 sg13g2_a22oi_1 _08928_ (.Y(_03373_),
    .B1(net3877),
    .B2(\jtag0.idr[16] ),
    .A2(net3887),
    .A1(\jtag0.idr[15] ));
 sg13g2_inv_1 _08929_ (.Y(_01269_),
    .A(_03373_));
 sg13g2_a22oi_1 _08930_ (.Y(_01268_),
    .B1(net3878),
    .B2(_01557_),
    .A2(net3888),
    .A1(_01558_));
 sg13g2_a22oi_1 _08931_ (.Y(_01267_),
    .B1(net3878),
    .B2(_01558_),
    .A2(net3888),
    .A1(_01559_));
 sg13g2_a22oi_1 _08932_ (.Y(_01266_),
    .B1(net3878),
    .B2(_01559_),
    .A2(net3888),
    .A1(_01560_));
 sg13g2_a22oi_1 _08933_ (.Y(_01265_),
    .B1(net3877),
    .B2(_01560_),
    .A2(net3887),
    .A1(_01561_));
 sg13g2_a22oi_1 _08934_ (.Y(_01264_),
    .B1(net3878),
    .B2(_01561_),
    .A2(net3888),
    .A1(_01562_));
 sg13g2_a22oi_1 _08935_ (.Y(_01263_),
    .B1(net3878),
    .B2(_01562_),
    .A2(net3888),
    .A1(_01563_));
 sg13g2_a22oi_1 _08936_ (.Y(_01262_),
    .B1(net3878),
    .B2(_01563_),
    .A2(net3888),
    .A1(_01564_));
 sg13g2_a22oi_1 _08937_ (.Y(_01261_),
    .B1(net3877),
    .B2(_01564_),
    .A2(net3887),
    .A1(_01565_));
 sg13g2_a22oi_1 _08938_ (.Y(_03374_),
    .B1(net3877),
    .B2(\jtag0.idr[7] ),
    .A2(net3887),
    .A1(\jtag0.idr[6] ));
 sg13g2_inv_1 _08939_ (.Y(_01260_),
    .A(_03374_));
 sg13g2_a22oi_1 _08940_ (.Y(_01259_),
    .B1(net3877),
    .B2(_01566_),
    .A2(net3887),
    .A1(_01567_));
 sg13g2_a22oi_1 _08941_ (.Y(_03375_),
    .B1(net3879),
    .B2(\jtag0.idr[5] ),
    .A2(net3889),
    .A1(\jtag0.idr[4] ));
 sg13g2_inv_1 _08942_ (.Y(_01258_),
    .A(_03375_));
 sg13g2_a22oi_1 _08943_ (.Y(_01257_),
    .B1(net3879),
    .B2(_01568_),
    .A2(net3889),
    .A1(_01569_));
 sg13g2_a22oi_1 _08944_ (.Y(_03376_),
    .B1(net3881),
    .B2(\jtag0.idr[3] ),
    .A2(net3891),
    .A1(\jtag0.idr[2] ));
 sg13g2_inv_1 _08945_ (.Y(_01256_),
    .A(_03376_));
 sg13g2_a22oi_1 _08946_ (.Y(_01255_),
    .B1(net3881),
    .B2(_01570_),
    .A2(net3891),
    .A1(_01571_));
 sg13g2_a22oi_1 _08947_ (.Y(_01254_),
    .B1(net3881),
    .B2(_01571_),
    .A2(net3891),
    .A1(_01572_));
 sg13g2_nand3_1 _08948_ (.B(\jtag0.ir[1] ),
    .C(\jtag0.ir[0] ),
    .A(\jtag0.ir[2] ),
    .Y(_03377_));
 sg13g2_mux2_1 _08949_ (.A0(\jtag0.stdi ),
    .A1(\jtag0.byp ),
    .S(_03377_),
    .X(_01253_));
 sg13g2_nand2_1 _08950_ (.Y(_03378_),
    .A(\jtag0.tapst[3] ),
    .B(net3926));
 sg13g2_nor2_2 _08951_ (.A(_01700_),
    .B(_02551_),
    .Y(_03379_));
 sg13g2_or2_1 _08952_ (.X(_03380_),
    .B(\jtag0.tapst[1] ),
    .A(net3927));
 sg13g2_nor2_1 _08953_ (.A(net3926),
    .B(_03380_),
    .Y(_03381_));
 sg13g2_a21oi_2 _08954_ (.B1(_03379_),
    .Y(_03382_),
    .A2(_03381_),
    .A1(_01700_));
 sg13g2_a22oi_1 _08955_ (.Y(_03383_),
    .B1(_03382_),
    .B2(\jtag0.ir[2] ),
    .A2(_03379_),
    .A1(\jtag0.irsh[2] ));
 sg13g2_inv_1 _08956_ (.Y(_01252_),
    .A(_03383_));
 sg13g2_a22oi_1 _08957_ (.Y(_03384_),
    .B1(_03382_),
    .B2(\jtag0.ir[1] ),
    .A2(_03379_),
    .A1(\jtag0.irsh[1] ));
 sg13g2_inv_1 _08958_ (.Y(_01251_),
    .A(_03384_));
 sg13g2_a22oi_1 _08959_ (.Y(_03385_),
    .B1(_03382_),
    .B2(\jtag0.ir[0] ),
    .A2(_03379_),
    .A1(\jtag0.irsh[0] ));
 sg13g2_inv_1 _08960_ (.Y(_01250_),
    .A(_03385_));
 sg13g2_and2_1 _08961_ (.A(net3050),
    .B(_02528_),
    .X(_03386_));
 sg13g2_nand2_2 _08962_ (.Y(_03387_),
    .A(net3050),
    .B(_02528_));
 sg13g2_nand2_1 _08963_ (.Y(_03388_),
    .A(_00580_),
    .B(net3048));
 sg13g2_o21ai_1 _08964_ (.B1(_03388_),
    .Y(_01113_),
    .A1(net3051),
    .A2(_02663_));
 sg13g2_nor2b_2 _08965_ (.A(_02528_),
    .B_N(net3050),
    .Y(_03389_));
 sg13g2_a22oi_1 _08966_ (.Y(_03390_),
    .B1(_03389_),
    .B2(_01747_),
    .A2(net3048),
    .A1(_00579_));
 sg13g2_o21ai_1 _08967_ (.B1(_03390_),
    .Y(_01112_),
    .A1(net3050),
    .A2(net3329));
 sg13g2_a22oi_1 _08968_ (.Y(_03391_),
    .B1(_03389_),
    .B2(_01746_),
    .A2(net3048),
    .A1(_00578_));
 sg13g2_o21ai_1 _08969_ (.B1(_03391_),
    .Y(_01111_),
    .A1(net3051),
    .A2(net3328));
 sg13g2_a22oi_1 _08970_ (.Y(_03392_),
    .B1(_03389_),
    .B2(_01745_),
    .A2(_03386_),
    .A1(_00577_));
 sg13g2_o21ai_1 _08971_ (.B1(_03392_),
    .Y(_01110_),
    .A1(net3051),
    .A2(_02927_));
 sg13g2_a22oi_1 _08972_ (.Y(_03393_),
    .B1(_03389_),
    .B2(_01744_),
    .A2(_03386_),
    .A1(_00576_));
 sg13g2_o21ai_1 _08973_ (.B1(_03393_),
    .Y(_01109_),
    .A1(net3051),
    .A2(net3327));
 sg13g2_a22oi_1 _08974_ (.Y(_03394_),
    .B1(_03389_),
    .B2(_01743_),
    .A2(net3048),
    .A1(_00575_));
 sg13g2_o21ai_1 _08975_ (.B1(_03394_),
    .Y(_01108_),
    .A1(net3051),
    .A2(net3326));
 sg13g2_a22oi_1 _08976_ (.Y(_03395_),
    .B1(_03389_),
    .B2(_01742_),
    .A2(net3048),
    .A1(_00574_));
 sg13g2_o21ai_1 _08977_ (.B1(_03395_),
    .Y(_01107_),
    .A1(_02469_),
    .A2(net3051));
 sg13g2_a22oi_1 _08978_ (.Y(_03396_),
    .B1(_03389_),
    .B2(_01741_),
    .A2(net3048),
    .A1(_00573_));
 sg13g2_o21ai_1 _08979_ (.B1(_03396_),
    .Y(_01106_),
    .A1(_02498_),
    .A2(net3051));
 sg13g2_a22oi_1 _08980_ (.Y(_01105_),
    .B1(_03389_),
    .B2(\uart0.txsh[1] ),
    .A2(net3048),
    .A1(_01574_));
 sg13g2_nor3_1 _08981_ (.A(\jtag0.ir[1] ),
    .B(\jtag0.ir[0] ),
    .C(_01705_),
    .Y(_03397_));
 sg13g2_a21oi_1 _08982_ (.A1(_01554_),
    .A2(_03377_),
    .Y(_03398_),
    .B1(_03397_));
 sg13g2_o21ai_1 _08983_ (.B1(_03398_),
    .Y(_03399_),
    .A1(\jtag0.byp ),
    .A2(_03377_));
 sg13g2_a21oi_1 _08984_ (.A1(\jtag0.idr[0] ),
    .A2(_03397_),
    .Y(_03400_),
    .B1(_01753_));
 sg13g2_a22oi_1 _08985_ (.Y(_03401_),
    .B1(_03399_),
    .B2(_03400_),
    .A2(_01753_),
    .A1(_01539_));
 sg13g2_nor2_1 _08986_ (.A(_03381_),
    .B(_03401_),
    .Y(_03402_));
 sg13g2_a21oi_1 _08987_ (.A1(_01706_),
    .A2(_03381_),
    .Y(pwmpin),
    .B1(_03402_));
 sg13g2_nand2b_1 _08988_ (.Y(_03403_),
    .B(net3925),
    .A_N(\ckd[2] ));
 sg13g2_and2_1 _08989_ (.A(net890),
    .B(_03403_),
    .X(_00000_));
 sg13g2_nor2b_1 _08990_ (.A(_02706_),
    .B_N(_03403_),
    .Y(_03404_));
 sg13g2_and2_1 _08991_ (.A(_02629_),
    .B(_03404_),
    .X(_00001_));
 sg13g2_nand2_1 _08992_ (.Y(_00002_),
    .A(_02711_),
    .B(_03403_));
 sg13g2_nand2_1 _08993_ (.Y(_03405_),
    .A(\pwmc[5] ),
    .B(\pwmc[7] ));
 sg13g2_nor3_2 _08994_ (.A(_00543_),
    .B(_00542_),
    .C(_03405_),
    .Y(_03406_));
 sg13g2_inv_1 _08995_ (.Y(_03407_),
    .A(_03406_));
 sg13g2_nor2_1 _08996_ (.A(\pwmc[0] ),
    .B(_03406_),
    .Y(_00004_));
 sg13g2_nand2_1 _08997_ (.Y(_03408_),
    .A(\pwmc[1] ),
    .B(\pwmc[0] ));
 sg13g2_nor2b_1 _08998_ (.A(_03406_),
    .B_N(_03408_),
    .Y(_03409_));
 sg13g2_o21ai_1 _08999_ (.B1(_03409_),
    .Y(_03410_),
    .A1(\pwmc[1] ),
    .A2(\pwmc[0] ));
 sg13g2_inv_1 _09000_ (.Y(_00005_),
    .A(_03410_));
 sg13g2_nor2_1 _09001_ (.A(_00542_),
    .B(_03409_),
    .Y(_03411_));
 sg13g2_a21oi_1 _09002_ (.A1(_00542_),
    .A2(_03408_),
    .Y(_00006_),
    .B1(_03411_));
 sg13g2_nand3_1 _09003_ (.B(\pwmc[0] ),
    .C(\pwmc[2] ),
    .A(\pwmc[1] ),
    .Y(_03412_));
 sg13g2_nor2_2 _09004_ (.A(_01703_),
    .B(_03412_),
    .Y(_03413_));
 sg13g2_and2_1 _09005_ (.A(_01703_),
    .B(_03412_),
    .X(_03414_));
 sg13g2_nor3_1 _09006_ (.A(_03406_),
    .B(_03413_),
    .C(_03414_),
    .Y(_00007_));
 sg13g2_nor3_1 _09007_ (.A(_00543_),
    .B(_03406_),
    .C(_03413_),
    .Y(_03415_));
 sg13g2_a21o_1 _09008_ (.A2(_03413_),
    .A1(_00543_),
    .B1(_03415_),
    .X(_00008_));
 sg13g2_a21oi_1 _09009_ (.A1(\pwmc[4] ),
    .A2(_03413_),
    .Y(_03416_),
    .B1(\pwmc[5] ));
 sg13g2_and3_1 _09010_ (.X(_03417_),
    .A(\pwmc[5] ),
    .B(\pwmc[4] ),
    .C(_03413_));
 sg13g2_nor3_1 _09011_ (.A(_03406_),
    .B(_03416_),
    .C(_03417_),
    .Y(_00009_));
 sg13g2_nand2_1 _09012_ (.Y(_03418_),
    .A(\pwmc[6] ),
    .B(_03417_));
 sg13g2_o21ai_1 _09013_ (.B1(_03407_),
    .Y(_03419_),
    .A1(\pwmc[6] ),
    .A2(_03417_));
 sg13g2_nor2b_1 _09014_ (.A(_03419_),
    .B_N(_03418_),
    .Y(_00010_));
 sg13g2_xor2_1 _09015_ (.B(_03418_),
    .A(\pwmc[7] ),
    .X(_03420_));
 sg13g2_nor2_1 _09016_ (.A(_03406_),
    .B(_03420_),
    .Y(_00011_));
 sg13g2_mux2_1 _09017_ (.A0(\cpu.PCreg0[18] ),
    .A1(\cpu.PCreg1[18] ),
    .S(net3633),
    .X(\cpu.PC[18] ));
 sg13g2_mux2_2 _09018_ (.A0(\cpu.PCreg0[19] ),
    .A1(\cpu.PCreg1[19] ),
    .S(net3632),
    .X(\cpu.PC[19] ));
 sg13g2_mux2_2 _09019_ (.A0(\cpu.PCreg0[20] ),
    .A1(\cpu.PCreg1[20] ),
    .S(net3631),
    .X(\cpu.PC[20] ));
 sg13g2_mux2_1 _09020_ (.A0(\cpu.PCreg0[21] ),
    .A1(\cpu.PCreg1[21] ),
    .S(net3632),
    .X(\cpu.PC[21] ));
 sg13g2_mux2_2 _09021_ (.A0(\cpu.PCreg0[22] ),
    .A1(\cpu.PCreg1[22] ),
    .S(net3632),
    .X(\cpu.PC[22] ));
 sg13g2_mux2_2 _09022_ (.A0(\cpu.PCreg0[23] ),
    .A1(\cpu.PCreg1[23] ),
    .S(net3632),
    .X(\cpu.PC[23] ));
 sg13g2_mux2_2 _09023_ (.A0(\cpu.PCreg0[24] ),
    .A1(\cpu.PCreg1[24] ),
    .S(net3632),
    .X(\cpu.PC[24] ));
 sg13g2_mux2_2 _09024_ (.A0(\cpu.PCreg0[25] ),
    .A1(\cpu.PCreg1[25] ),
    .S(net3632),
    .X(\cpu.PC[25] ));
 sg13g2_mux2_2 _09025_ (.A0(\cpu.PCreg0[26] ),
    .A1(\cpu.PCreg1[26] ),
    .S(net3633),
    .X(\cpu.PC[26] ));
 sg13g2_mux2_2 _09026_ (.A0(\cpu.PCreg0[27] ),
    .A1(\cpu.PCreg1[27] ),
    .S(net3634),
    .X(\cpu.PC[27] ));
 sg13g2_mux2_2 _09027_ (.A0(\cpu.PCreg0[28] ),
    .A1(\cpu.PCreg1[28] ),
    .S(net3633),
    .X(\cpu.PC[28] ));
 sg13g2_and2_2 _09028_ (.A(_02419_),
    .B(net3142),
    .X(_03421_));
 sg13g2_nor2_2 _09029_ (.A(_02414_),
    .B(_02418_),
    .Y(_03422_));
 sg13g2_nand2_1 _09030_ (.Y(_03423_),
    .A(_03345_),
    .B(_03422_));
 sg13g2_nand2_1 _09031_ (.Y(_03424_),
    .A(net3122),
    .B(net3128));
 sg13g2_nor2b_2 _09032_ (.A(_03424_),
    .B_N(_02408_),
    .Y(_03425_));
 sg13g2_nor2_2 _09033_ (.A(_02408_),
    .B(_03424_),
    .Y(_03426_));
 sg13g2_inv_1 _09034_ (.Y(_03427_),
    .A(_03426_));
 sg13g2_a22oi_1 _09035_ (.Y(_03428_),
    .B1(_03426_),
    .B2(\tcount[0] ),
    .A2(_03425_),
    .A1(\irqen[0] ));
 sg13g2_nand2_1 _09036_ (.Y(_03429_),
    .A(_03423_),
    .B(_03428_));
 sg13g2_a221oi_1 _09037_ (.B2(\uart0.rxvalid ),
    .C1(_03429_),
    .B1(_03421_),
    .A1(\uart0.q[0] ),
    .Y(_03430_),
    .A2(net3117));
 sg13g2_nand2b_1 _09038_ (.Y(_03431_),
    .B(net3098),
    .A_N(_03430_));
 sg13g2_nand4_1 _09039_ (.B(_02395_),
    .C(_02398_),
    .A(_02390_),
    .Y(_03432_),
    .D(_02400_));
 sg13g2_nor3_2 _09040_ (.A(_01767_),
    .B(_02387_),
    .C(_03432_),
    .Y(_03433_));
 sg13g2_or3_2 _09041_ (.A(_01767_),
    .B(_02387_),
    .C(_03432_),
    .X(_03434_));
 sg13g2_a21oi_1 _09042_ (.A1(\xdi[0] ),
    .A2(net3096),
    .Y(_03435_),
    .B1(net3091));
 sg13g2_nand2_1 _09043_ (.Y(\cdi[0] ),
    .A(_03431_),
    .B(_03435_));
 sg13g2_nor4_1 _09044_ (.A(_02388_),
    .B(_02389_),
    .C(_02403_),
    .D(_03427_),
    .Y(_03436_));
 sg13g2_and2_1 _09045_ (.A(\tcount[16] ),
    .B(net3086),
    .X(_03437_));
 sg13g2_nand2_1 _09046_ (.Y(_03438_),
    .A(net3126),
    .B(_03223_));
 sg13g2_and2_1 _09047_ (.A(net3141),
    .B(_03149_),
    .X(_03439_));
 sg13g2_inv_1 _09048_ (.Y(_03440_),
    .A(_03439_));
 sg13g2_nor2_2 _09049_ (.A(net3126),
    .B(_03439_),
    .Y(_03441_));
 sg13g2_nand2_2 _09050_ (.Y(_03442_),
    .A(net3142),
    .B(_03224_));
 sg13g2_nand2b_2 _09051_ (.Y(_03443_),
    .B(_03223_),
    .A_N(net3141));
 sg13g2_or2_1 _09052_ (.X(_03444_),
    .B(_03223_),
    .A(net3141));
 sg13g2_nand2_2 _09053_ (.Y(_03445_),
    .A(net3141),
    .B(_03223_));
 sg13g2_nand2_2 _09054_ (.Y(_03446_),
    .A(_03444_),
    .B(_03445_));
 sg13g2_nand2_1 _09055_ (.Y(_03447_),
    .A(_03441_),
    .B(_03446_));
 sg13g2_nand3_1 _09056_ (.B(_03438_),
    .C(_03447_),
    .A(net3122),
    .Y(_03448_));
 sg13g2_nor2_1 _09057_ (.A(net3121),
    .B(_03150_),
    .Y(_03449_));
 sg13g2_a21o_1 _09058_ (.A2(_03449_),
    .A1(_03444_),
    .B1(net3122),
    .X(_03450_));
 sg13g2_nor2_1 _09059_ (.A(net3125),
    .B(_03444_),
    .Y(_03451_));
 sg13g2_inv_2 _09060_ (.Y(_03452_),
    .A(_03451_));
 sg13g2_nor2_1 _09061_ (.A(net3141),
    .B(net3124),
    .Y(_03453_));
 sg13g2_nand2b_1 _09062_ (.Y(_03454_),
    .B(_03149_),
    .A_N(net3142));
 sg13g2_a21oi_1 _09063_ (.A1(_03223_),
    .A2(_03453_),
    .Y(_03455_),
    .B1(net3126));
 sg13g2_and2_1 _09064_ (.A(_03452_),
    .B(_03455_),
    .X(_03456_));
 sg13g2_o21ai_1 _09065_ (.B1(_03448_),
    .Y(_03457_),
    .A1(_03450_),
    .A2(_03456_));
 sg13g2_a221oi_1 _09066_ (.B2(_03457_),
    .C1(_03437_),
    .B1(net3091),
    .A1(\xdi[16] ),
    .Y(_03458_),
    .A2(net3092));
 sg13g2_inv_1 _09067_ (.Y(\cdi[16] ),
    .A(_03458_));
 sg13g2_nand2_1 _09068_ (.Y(_03459_),
    .A(_03341_),
    .B(_03422_));
 sg13g2_a22oi_1 _09069_ (.Y(_03460_),
    .B1(_03426_),
    .B2(\tcount[1] ),
    .A2(_03425_),
    .A1(\irqen[1] ));
 sg13g2_a22oi_1 _09070_ (.Y(_03461_),
    .B1(_02425_),
    .B2(_03421_),
    .A2(net3117),
    .A1(\uart0.q[1] ));
 sg13g2_nand3_1 _09071_ (.B(_03460_),
    .C(_03461_),
    .A(_03459_),
    .Y(_03462_));
 sg13g2_a21oi_1 _09072_ (.A1(net3099),
    .A2(_03462_),
    .Y(_03463_),
    .B1(net3091));
 sg13g2_o21ai_1 _09073_ (.B1(_03463_),
    .Y(\cdi[1] ),
    .A1(_01734_),
    .A2(_02570_));
 sg13g2_nand2_1 _09074_ (.Y(_03464_),
    .A(net3127),
    .B(_03446_));
 sg13g2_a21o_1 _09075_ (.A2(_03454_),
    .A1(_03442_),
    .B1(net3127),
    .X(_03465_));
 sg13g2_nand3_1 _09076_ (.B(_03464_),
    .C(_03465_),
    .A(net3122),
    .Y(_03466_));
 sg13g2_nor2_1 _09077_ (.A(_03439_),
    .B(_03451_),
    .Y(_03467_));
 sg13g2_o21ai_1 _09078_ (.B1(net3119),
    .Y(_03468_),
    .A1(net3120),
    .A2(_03467_));
 sg13g2_nor2_2 _09079_ (.A(net3125),
    .B(_03443_),
    .Y(_03469_));
 sg13g2_nand2_1 _09080_ (.Y(_03470_),
    .A(net3120),
    .B(_03224_));
 sg13g2_nor2b_2 _09081_ (.A(_03441_),
    .B_N(_03470_),
    .Y(_03471_));
 sg13g2_inv_1 _09082_ (.Y(_03472_),
    .A(_03471_));
 sg13g2_nor2_1 _09083_ (.A(_03469_),
    .B(_03471_),
    .Y(_03473_));
 sg13g2_o21ai_1 _09084_ (.B1(_03466_),
    .Y(_03474_),
    .A1(_03468_),
    .A2(_03473_));
 sg13g2_and2_1 _09085_ (.A(\xdi[17] ),
    .B(net3094),
    .X(_03475_));
 sg13g2_a221oi_1 _09086_ (.B2(net3090),
    .C1(_03475_),
    .B1(_03474_),
    .A1(\tcount[17] ),
    .Y(_03476_),
    .A2(net3086));
 sg13g2_inv_1 _09087_ (.Y(\cdi[17] ),
    .A(_03476_));
 sg13g2_nor2_1 _09088_ (.A(net3120),
    .B(_03440_),
    .Y(_03477_));
 sg13g2_o21ai_1 _09089_ (.B1(net3118),
    .Y(_03478_),
    .A1(net3120),
    .A2(_03440_));
 sg13g2_nor2_2 _09090_ (.A(net3124),
    .B(_03223_),
    .Y(_03479_));
 sg13g2_or2_1 _09091_ (.X(_03480_),
    .B(_03479_),
    .A(net3141));
 sg13g2_a21oi_1 _09092_ (.A1(_03441_),
    .A2(_03480_),
    .Y(_03481_),
    .B1(_03478_));
 sg13g2_nor2_1 _09093_ (.A(net3121),
    .B(_03445_),
    .Y(_03482_));
 sg13g2_nor2_1 _09094_ (.A(_03454_),
    .B(_03470_),
    .Y(_03483_));
 sg13g2_nor3_1 _09095_ (.A(net3118),
    .B(_03482_),
    .C(_03483_),
    .Y(_03484_));
 sg13g2_nand2b_1 _09096_ (.Y(_03485_),
    .B(_03433_),
    .A_N(_03484_));
 sg13g2_nand2_1 _09097_ (.Y(_03486_),
    .A(\uart0.q[2] ),
    .B(net3117));
 sg13g2_nand2b_1 _09098_ (.Y(_03487_),
    .B(_03421_),
    .A_N(\uart0.urxbuffer[8] ));
 sg13g2_nand2_1 _09099_ (.Y(_03488_),
    .A(\irqen[2] ),
    .B(_03425_));
 sg13g2_a22oi_1 _09100_ (.Y(_03489_),
    .B1(_03426_),
    .B2(\tcount[2] ),
    .A2(_03422_),
    .A1(_03337_));
 sg13g2_nand4_1 _09101_ (.B(_03487_),
    .C(_03488_),
    .A(_03486_),
    .Y(_03490_),
    .D(_03489_));
 sg13g2_a22oi_1 _09102_ (.Y(_03491_),
    .B1(_03490_),
    .B2(net3099),
    .A2(net3094),
    .A1(\xdi[2] ));
 sg13g2_o21ai_1 _09103_ (.B1(_03491_),
    .Y(\cdi[2] ),
    .A1(_03481_),
    .A2(_03485_));
 sg13g2_nor4_1 _09104_ (.A(net3119),
    .B(_03434_),
    .C(_03454_),
    .D(_03470_),
    .Y(_03492_));
 sg13g2_a221oi_1 _09105_ (.B2(\tcount[18] ),
    .C1(_03492_),
    .B1(net3087),
    .A1(\xdi[18] ),
    .Y(_03493_),
    .A2(net3093));
 sg13g2_inv_1 _09106_ (.Y(\cdi[18] ),
    .A(_03493_));
 sg13g2_nand2_1 _09107_ (.Y(_03494_),
    .A(_03333_),
    .B(_03422_));
 sg13g2_a22oi_1 _09108_ (.Y(_03495_),
    .B1(_03426_),
    .B2(\tcount[3] ),
    .A2(_03425_),
    .A1(\irqen[3] ));
 sg13g2_a22oi_1 _09109_ (.Y(_03496_),
    .B1(_03421_),
    .B2(\uart0.rxoverr ),
    .A2(net3117),
    .A1(\uart0.q[3] ));
 sg13g2_nand3_1 _09110_ (.B(_03495_),
    .C(_03496_),
    .A(_03494_),
    .Y(_03497_));
 sg13g2_a21oi_1 _09111_ (.A1(net3141),
    .A2(net3124),
    .Y(_03498_),
    .B1(net3126));
 sg13g2_a21oi_1 _09112_ (.A1(net3127),
    .A2(_03440_),
    .Y(_03499_),
    .B1(net3123));
 sg13g2_nand2b_1 _09113_ (.Y(_03500_),
    .B(_03499_),
    .A_N(_03498_));
 sg13g2_a22oi_1 _09114_ (.Y(_03501_),
    .B1(_03497_),
    .B2(net3098),
    .A2(net3092),
    .A1(\xdi[3] ));
 sg13g2_o21ai_1 _09115_ (.B1(_03501_),
    .Y(\cdi[3] ),
    .A1(_03434_),
    .A2(_03500_));
 sg13g2_a22oi_1 _09116_ (.Y(_03502_),
    .B1(net3086),
    .B2(\tcount[19] ),
    .A2(net3092),
    .A1(\xdi[19] ));
 sg13g2_inv_1 _09117_ (.Y(\cdi[19] ),
    .A(_03502_));
 sg13g2_nor4_1 _09118_ (.A(_01540_),
    .B(\uart0.q[7] ),
    .C(\uart0.q[6] ),
    .D(\uart0.q[3] ),
    .Y(_03503_));
 sg13g2_nand4_1 _09119_ (.B(\uart0.q[1] ),
    .C(\uart0.q[0] ),
    .A(_01541_),
    .Y(_03504_),
    .D(_03503_));
 sg13g2_nor3_2 _09120_ (.A(\uart0.q[5] ),
    .B(\uart0.q[4] ),
    .C(_03504_),
    .Y(_03505_));
 sg13g2_a22oi_1 _09121_ (.Y(_03506_),
    .B1(_03505_),
    .B2(_03421_),
    .A2(_03426_),
    .A1(\tcount[4] ));
 sg13g2_inv_1 _09122_ (.Y(_03507_),
    .A(_03506_));
 sg13g2_a221oi_1 _09123_ (.B2(\irqen[4] ),
    .C1(_03507_),
    .B1(_03425_),
    .A1(\uart0.q[4] ),
    .Y(_03508_),
    .A2(net3117));
 sg13g2_nand2b_1 _09124_ (.Y(_03509_),
    .B(net3098),
    .A_N(_03508_));
 sg13g2_nor3_1 _09125_ (.A(_03449_),
    .B(_03469_),
    .C(_03479_),
    .Y(_03510_));
 sg13g2_o21ai_1 _09126_ (.B1(_03466_),
    .Y(_03511_),
    .A1(_03478_),
    .A2(_03510_));
 sg13g2_a22oi_1 _09127_ (.Y(_03512_),
    .B1(net3090),
    .B2(_03511_),
    .A2(net3093),
    .A1(\xdi[4] ));
 sg13g2_nand2_2 _09128_ (.Y(\cdi[4] ),
    .A(_03509_),
    .B(_03512_));
 sg13g2_nor2_1 _09129_ (.A(_03451_),
    .B(_03471_),
    .Y(_03513_));
 sg13g2_nor2_1 _09130_ (.A(net3125),
    .B(_03464_),
    .Y(_03514_));
 sg13g2_nor4_1 _09131_ (.A(_03434_),
    .B(_03450_),
    .C(_03513_),
    .D(_03514_),
    .Y(_03515_));
 sg13g2_a221oi_1 _09132_ (.B2(\tcount[20] ),
    .C1(_03515_),
    .B1(net3086),
    .A1(\xdi[20] ),
    .Y(_03516_),
    .A2(net3093));
 sg13g2_inv_1 _09133_ (.Y(\cdi[20] ),
    .A(_03516_));
 sg13g2_nand2_1 _09134_ (.Y(_03517_),
    .A(udirty),
    .B(_03421_));
 sg13g2_nand2b_1 _09135_ (.Y(_03518_),
    .B(net3126),
    .A_N(net3141));
 sg13g2_nand2b_1 _09136_ (.Y(_03519_),
    .B(_03498_),
    .A_N(_03446_));
 sg13g2_o21ai_1 _09137_ (.B1(_03519_),
    .Y(_03520_),
    .A1(_03479_),
    .A2(_03518_));
 sg13g2_nand2_1 _09138_ (.Y(_03521_),
    .A(net3091),
    .B(_03448_));
 sg13g2_a21oi_1 _09139_ (.A1(net3118),
    .A2(_03520_),
    .Y(_03522_),
    .B1(_03521_));
 sg13g2_a22oi_1 _09140_ (.Y(_03523_),
    .B1(_03426_),
    .B2(\tcount[5] ),
    .A2(net3117),
    .A1(\uart0.q[5] ));
 sg13g2_nand2_1 _09141_ (.Y(_03524_),
    .A(_03517_),
    .B(_03523_));
 sg13g2_a221oi_1 _09142_ (.B2(net3099),
    .C1(_03522_),
    .B1(_03524_),
    .A1(\xdi[5] ),
    .Y(_03525_),
    .A2(net3092));
 sg13g2_inv_1 _09143_ (.Y(\cdi[5] ),
    .A(_03525_));
 sg13g2_nand2_1 _09144_ (.Y(_03526_),
    .A(net3127),
    .B(_03443_));
 sg13g2_a21o_1 _09145_ (.A2(_03446_),
    .A1(net3124),
    .B1(net3126),
    .X(_03527_));
 sg13g2_and4_2 _09146_ (.A(net3123),
    .B(net3090),
    .C(_03526_),
    .D(_03527_),
    .X(_03528_));
 sg13g2_a221oi_1 _09147_ (.B2(\tcount[21] ),
    .C1(_03528_),
    .B1(net3089),
    .A1(\xdi[21] ),
    .Y(_03529_),
    .A2(net3093));
 sg13g2_inv_1 _09148_ (.Y(\cdi[21] ),
    .A(_03529_));
 sg13g2_nor2_1 _09149_ (.A(net3125),
    .B(_03445_),
    .Y(_03530_));
 sg13g2_nor2_2 _09150_ (.A(net3120),
    .B(_03530_),
    .Y(_03531_));
 sg13g2_inv_1 _09151_ (.Y(_03532_),
    .A(_03531_));
 sg13g2_nand2_1 _09152_ (.Y(_03533_),
    .A(_03445_),
    .B(_03498_));
 sg13g2_a21oi_1 _09153_ (.A1(_03532_),
    .A2(_03533_),
    .Y(_03534_),
    .B1(_03478_));
 sg13g2_nand2_1 _09154_ (.Y(_03535_),
    .A(pwmirq),
    .B(_03421_));
 sg13g2_a22oi_1 _09155_ (.Y(_03536_),
    .B1(_03426_),
    .B2(\tcount[6] ),
    .A2(net3117),
    .A1(\uart0.q[6] ));
 sg13g2_nand2_1 _09156_ (.Y(_03537_),
    .A(_03535_),
    .B(_03536_));
 sg13g2_a22oi_1 _09157_ (.Y(_03538_),
    .B1(_03537_),
    .B2(net3099),
    .A2(net3096),
    .A1(\xdi[6] ));
 sg13g2_o21ai_1 _09158_ (.B1(_03538_),
    .Y(\cdi[6] ),
    .A1(_03485_),
    .A2(_03534_));
 sg13g2_a21oi_2 _09159_ (.B1(_03528_),
    .Y(_03539_),
    .A2(net3093),
    .A1(\xdi[22] ));
 sg13g2_nand2_1 _09160_ (.Y(_03540_),
    .A(net3126),
    .B(_03224_));
 sg13g2_a21oi_1 _09161_ (.A1(_03467_),
    .A2(_03540_),
    .Y(_03541_),
    .B1(_03468_));
 sg13g2_a22oi_1 _09162_ (.Y(_03542_),
    .B1(_03541_),
    .B2(net3090),
    .A2(net3086),
    .A1(\tcount[22] ));
 sg13g2_nand2_2 _09163_ (.Y(\cdi[22] ),
    .A(_03539_),
    .B(_03542_));
 sg13g2_nand3_1 _09164_ (.B(net3098),
    .C(net3117),
    .A(\uart0.q[7] ),
    .Y(_03543_));
 sg13g2_nand2_1 _09165_ (.Y(_03544_),
    .A(\tcount[7] ),
    .B(net3088));
 sg13g2_a21o_1 _09166_ (.A2(_03479_),
    .A1(net3142),
    .B1(_03530_),
    .X(_03545_));
 sg13g2_nand2_1 _09167_ (.Y(_03546_),
    .A(net3121),
    .B(_03452_));
 sg13g2_o21ai_1 _09168_ (.B1(_03526_),
    .Y(_03547_),
    .A1(_03545_),
    .A2(_03546_));
 sg13g2_and2_1 _09169_ (.A(net3125),
    .B(_03446_),
    .X(_03548_));
 sg13g2_nor2_1 _09170_ (.A(_03149_),
    .B(_03442_),
    .Y(_03549_));
 sg13g2_nor2_1 _09171_ (.A(_03548_),
    .B(_03549_),
    .Y(_03550_));
 sg13g2_o21ai_1 _09172_ (.B1(net3120),
    .Y(_03551_),
    .A1(_03548_),
    .A2(_03549_));
 sg13g2_a21oi_1 _09173_ (.A1(_03470_),
    .A2(_03550_),
    .Y(_03552_),
    .B1(net3123));
 sg13g2_a22oi_1 _09174_ (.Y(_03553_),
    .B1(_03551_),
    .B2(_03552_),
    .A2(_03547_),
    .A1(net3123));
 sg13g2_a22oi_1 _09175_ (.Y(_03554_),
    .B1(net3091),
    .B2(_03553_),
    .A2(net3092),
    .A1(\xdi[7] ));
 sg13g2_nand3_1 _09176_ (.B(_03544_),
    .C(_03554_),
    .A(_03543_),
    .Y(\cdi[7] ));
 sg13g2_nand2_1 _09177_ (.Y(_03555_),
    .A(net3118),
    .B(net3090));
 sg13g2_nor2_1 _09178_ (.A(_03531_),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_and4_1 _09179_ (.A(net3119),
    .B(net3090),
    .C(_03532_),
    .D(_03545_),
    .X(_03557_));
 sg13g2_nand3_1 _09180_ (.B(_03438_),
    .C(_03518_),
    .A(net3122),
    .Y(_03558_));
 sg13g2_nor2_1 _09181_ (.A(_03472_),
    .B(_03558_),
    .Y(_03559_));
 sg13g2_inv_1 _09182_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_nor4_1 _09183_ (.A(_01767_),
    .B(_02387_),
    .C(_03432_),
    .D(_03560_),
    .Y(_03561_));
 sg13g2_a221oi_1 _09184_ (.B2(\tcount[23] ),
    .C1(_03561_),
    .B1(net3089),
    .A1(\xdi[23] ),
    .Y(_03562_),
    .A2(net3093));
 sg13g2_nand2b_2 _09185_ (.Y(\cdi[23] ),
    .B(_03562_),
    .A_N(_03557_));
 sg13g2_o21ai_1 _09186_ (.B1(_03540_),
    .Y(_03563_),
    .A1(_03479_),
    .A2(_03527_));
 sg13g2_nand2_1 _09187_ (.Y(_03564_),
    .A(net3122),
    .B(_03563_));
 sg13g2_o21ai_1 _09188_ (.B1(net3118),
    .Y(_03565_),
    .A1(_03469_),
    .A2(_03483_));
 sg13g2_a21oi_1 _09189_ (.A1(_03564_),
    .A2(_03565_),
    .Y(_03566_),
    .B1(_03434_));
 sg13g2_a221oi_1 _09190_ (.B2(\tcount[8] ),
    .C1(_03566_),
    .B1(net3088),
    .A1(\xdi[8] ),
    .Y(_03567_),
    .A2(net3094));
 sg13g2_inv_1 _09191_ (.Y(\cdi[8] ),
    .A(_03567_));
 sg13g2_and2_1 _09192_ (.A(net3092),
    .B(_03329_),
    .X(_03568_));
 sg13g2_nor2_1 _09193_ (.A(net3127),
    .B(_03469_),
    .Y(_03569_));
 sg13g2_nor2b_1 _09194_ (.A(net3122),
    .B_N(_03540_),
    .Y(_03570_));
 sg13g2_o21ai_1 _09195_ (.B1(_03570_),
    .Y(_03571_),
    .A1(_03477_),
    .A2(_03549_));
 sg13g2_o21ai_1 _09196_ (.B1(_03571_),
    .Y(_03572_),
    .A1(_03558_),
    .A2(_03569_));
 sg13g2_a221oi_1 _09197_ (.B2(net3090),
    .C1(_03568_),
    .B1(_03572_),
    .A1(\tcount[24] ),
    .Y(_03573_),
    .A2(net3086));
 sg13g2_inv_1 _09198_ (.Y(\cdi[24] ),
    .A(_03573_));
 sg13g2_a21oi_1 _09199_ (.A1(net3124),
    .A2(_03442_),
    .Y(_03574_),
    .B1(net3120));
 sg13g2_a21o_1 _09200_ (.A2(_03443_),
    .A1(_03441_),
    .B1(_03574_),
    .X(_03575_));
 sg13g2_a22oi_1 _09201_ (.Y(_03576_),
    .B1(net3091),
    .B2(_03484_),
    .A2(net3094),
    .A1(\xdi[9] ));
 sg13g2_o21ai_1 _09202_ (.B1(_03576_),
    .Y(_03577_),
    .A1(_03555_),
    .A2(_03575_));
 sg13g2_a21o_2 _09203_ (.A2(net3087),
    .A1(\tcount[9] ),
    .B1(_03577_),
    .X(\cdi[9] ));
 sg13g2_o21ai_1 _09204_ (.B1(_03531_),
    .Y(_03578_),
    .A1(net3124),
    .A2(_03442_));
 sg13g2_nand2_1 _09205_ (.Y(_03579_),
    .A(_03533_),
    .B(_03578_));
 sg13g2_a22oi_1 _09206_ (.Y(_03580_),
    .B1(net3087),
    .B2(\tcount[25] ),
    .A2(_03325_),
    .A1(net3095));
 sg13g2_o21ai_1 _09207_ (.B1(_03580_),
    .Y(\cdi[25] ),
    .A1(_03555_),
    .A2(_03579_));
 sg13g2_inv_1 _09208_ (.Y(_03581_),
    .A(\cdi[25] ));
 sg13g2_o21ai_1 _09209_ (.B1(_03471_),
    .Y(_03582_),
    .A1(net3120),
    .A2(_03453_));
 sg13g2_a22oi_1 _09210_ (.Y(_03583_),
    .B1(net3087),
    .B2(\tcount[10] ),
    .A2(net3095),
    .A1(\xdi[10] ));
 sg13g2_o21ai_1 _09211_ (.B1(_03583_),
    .Y(\cdi[10] ),
    .A1(_03555_),
    .A2(_03582_));
 sg13g2_nand2b_1 _09212_ (.Y(_03584_),
    .B(_03556_),
    .A_N(_03441_));
 sg13g2_a22oi_1 _09213_ (.Y(_03585_),
    .B1(net3087),
    .B2(\tcount[26] ),
    .A2(_03321_),
    .A1(net3095));
 sg13g2_nand2_2 _09214_ (.Y(\cdi[26] ),
    .A(_03584_),
    .B(_03585_));
 sg13g2_nand2_2 _09215_ (.Y(_03586_),
    .A(_03471_),
    .B(_03556_));
 sg13g2_a22oi_1 _09216_ (.Y(_03587_),
    .B1(net3088),
    .B2(\tcount[11] ),
    .A2(net3096),
    .A1(\xdi[11] ));
 sg13g2_nand2_2 _09217_ (.Y(\cdi[11] ),
    .A(_03586_),
    .B(_03587_));
 sg13g2_inv_1 _09218_ (.Y(_03588_),
    .A(\cdi[11] ));
 sg13g2_a22oi_1 _09219_ (.Y(_03589_),
    .B1(net3087),
    .B2(\tcount[27] ),
    .A2(_03317_),
    .A1(net3095));
 sg13g2_nand2_2 _09220_ (.Y(\cdi[27] ),
    .A(_03586_),
    .B(_03589_));
 sg13g2_nand2_1 _09221_ (.Y(_03590_),
    .A(\tcount[12] ),
    .B(net3088));
 sg13g2_nor2_2 _09222_ (.A(_03473_),
    .B(_03558_),
    .Y(_03591_));
 sg13g2_a22oi_1 _09223_ (.Y(_03592_),
    .B1(net3090),
    .B2(_03591_),
    .A2(net3094),
    .A1(\xdi[12] ));
 sg13g2_and3_1 _09224_ (.X(_03593_),
    .A(_03586_),
    .B(_03590_),
    .C(_03592_));
 sg13g2_inv_1 _09225_ (.Y(\cdi[12] ),
    .A(_03593_));
 sg13g2_a22oi_1 _09226_ (.Y(_03594_),
    .B1(net3087),
    .B2(\tcount[28] ),
    .A2(_03314_),
    .A1(net3094));
 sg13g2_and2_2 _09227_ (.A(_03586_),
    .B(_03594_),
    .X(_03595_));
 sg13g2_inv_1 _09228_ (.Y(\cdi[28] ),
    .A(_03595_));
 sg13g2_a221oi_1 _09229_ (.B2(\tcount[13] ),
    .C1(_03528_),
    .B1(net3089),
    .A1(\xdi[13] ),
    .Y(_03596_),
    .A2(net3093));
 sg13g2_inv_1 _09230_ (.Y(\cdi[13] ),
    .A(_03596_));
 sg13g2_nor2_1 _09231_ (.A(net3127),
    .B(_03548_),
    .Y(_03597_));
 sg13g2_nor4_2 _09232_ (.A(net3123),
    .B(_03434_),
    .C(_03531_),
    .Y(_03598_),
    .D(_03597_));
 sg13g2_a221oi_1 _09233_ (.B2(\tcount[29] ),
    .C1(_03598_),
    .B1(net3088),
    .A1(net3094),
    .Y(_03599_),
    .A2(_03308_));
 sg13g2_inv_1 _09234_ (.Y(\cdi[29] ),
    .A(_03599_));
 sg13g2_nand2b_1 _09235_ (.Y(_03600_),
    .B(_03597_),
    .A_N(_03469_));
 sg13g2_a21oi_1 _09236_ (.A1(net3126),
    .A2(_03452_),
    .Y(_03601_),
    .B1(_03455_));
 sg13g2_a21oi_1 _09237_ (.A1(_03518_),
    .A2(_03600_),
    .Y(_03602_),
    .B1(net3118));
 sg13g2_a21oi_1 _09238_ (.A1(net3118),
    .A2(_03601_),
    .Y(_03603_),
    .B1(_03602_));
 sg13g2_nor2_1 _09239_ (.A(_03434_),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_a221oi_1 _09240_ (.B2(\tcount[14] ),
    .C1(_03604_),
    .B1(net3086),
    .A1(\xdi[14] ),
    .Y(_03605_),
    .A2(net3092));
 sg13g2_inv_1 _09241_ (.Y(\cdi[14] ),
    .A(_03605_));
 sg13g2_a221oi_1 _09242_ (.B2(\tcount[30] ),
    .C1(_03598_),
    .B1(net3088),
    .A1(net3094),
    .Y(_03606_),
    .A2(_03302_));
 sg13g2_inv_2 _09243_ (.Y(\cdi[30] ),
    .A(_03606_));
 sg13g2_a21oi_1 _09244_ (.A1(_03480_),
    .A2(_03499_),
    .Y(_03607_),
    .B1(_03591_));
 sg13g2_and2_1 _09245_ (.A(net3091),
    .B(_03607_),
    .X(_03608_));
 sg13g2_a221oi_1 _09246_ (.B2(\tcount[15] ),
    .C1(_03608_),
    .B1(net3086),
    .A1(\xdi[15] ),
    .Y(_03609_),
    .A2(net3092));
 sg13g2_inv_1 _09247_ (.Y(\cdi[15] ),
    .A(_03609_));
 sg13g2_a22oi_1 _09248_ (.Y(_03610_),
    .B1(net3087),
    .B2(\tcount[31] ),
    .A2(_03299_),
    .A1(net3095));
 sg13g2_nor2b_2 _09249_ (.A(_03598_),
    .B_N(_03610_),
    .Y(_03611_));
 sg13g2_inv_1 _09250_ (.Y(\cdi[31] ),
    .A(_03611_));
 sg13g2_nor2_1 _09251_ (.A(\uart0.txdiv[0] ),
    .B(_03387_),
    .Y(_00021_));
 sg13g2_xnor2_1 _09252_ (.Y(_03612_),
    .A(\uart0.txdiv[0] ),
    .B(\uart0.txdiv[1] ));
 sg13g2_nor2_1 _09253_ (.A(_03387_),
    .B(_03612_),
    .Y(_00022_));
 sg13g2_and3_1 _09254_ (.X(_03613_),
    .A(\uart0.txdiv[0] ),
    .B(\uart0.txdiv[1] ),
    .C(\uart0.txdiv[2] ));
 sg13g2_a21oi_1 _09255_ (.A1(\uart0.txdiv[0] ),
    .A2(\uart0.txdiv[1] ),
    .Y(_03614_),
    .B1(\uart0.txdiv[2] ));
 sg13g2_nor3_1 _09256_ (.A(_03387_),
    .B(_03613_),
    .C(_03614_),
    .Y(_00023_));
 sg13g2_and2_1 _09257_ (.A(\uart0.txdiv[3] ),
    .B(_03613_),
    .X(_03615_));
 sg13g2_nor2_1 _09258_ (.A(\uart0.txdiv[3] ),
    .B(_03613_),
    .Y(_03616_));
 sg13g2_nor3_1 _09259_ (.A(_03387_),
    .B(_03615_),
    .C(_03616_),
    .Y(_00024_));
 sg13g2_nand2_1 _09260_ (.Y(_03617_),
    .A(\uart0.txdiv[4] ),
    .B(_03615_));
 sg13g2_o21ai_1 _09261_ (.B1(net3048),
    .Y(_03618_),
    .A1(\uart0.txdiv[4] ),
    .A2(_03615_));
 sg13g2_nor2b_1 _09262_ (.A(_03618_),
    .B_N(_03617_),
    .Y(_00025_));
 sg13g2_xor2_1 _09263_ (.B(_03617_),
    .A(\uart0.txdiv[5] ),
    .X(_03619_));
 sg13g2_nor2_1 _09264_ (.A(_03387_),
    .B(_03619_),
    .Y(_00026_));
 sg13g2_xor2_1 _09265_ (.B(\uart0.rxreg[1] ),
    .A(\uart0.rxreg[0] ),
    .X(_03620_));
 sg13g2_nand3b_1 _09266_ (.B(\uart0.rxdiv[1] ),
    .C(\uart0.rxdiv[5] ),
    .Y(_03621_),
    .A_N(\uart0.rxdiv[0] ));
 sg13g2_nor4_1 _09267_ (.A(\uart0.rxdiv[3] ),
    .B(\uart0.rxdiv[2] ),
    .C(\uart0.rxdiv[4] ),
    .D(_03621_),
    .Y(_03622_));
 sg13g2_or2_2 _09268_ (.X(_03623_),
    .B(_03622_),
    .A(_03620_));
 sg13g2_nor2_1 _09269_ (.A(\uart0.rxdiv[0] ),
    .B(_03623_),
    .Y(_00015_));
 sg13g2_and2_1 _09270_ (.A(\uart0.rxdiv[0] ),
    .B(\uart0.rxdiv[1] ),
    .X(_03624_));
 sg13g2_nor3_1 _09271_ (.A(_02536_),
    .B(_03623_),
    .C(_03624_),
    .Y(_00016_));
 sg13g2_nor2_1 _09272_ (.A(\uart0.rxdiv[2] ),
    .B(_03624_),
    .Y(_03625_));
 sg13g2_and2_1 _09273_ (.A(\uart0.rxdiv[2] ),
    .B(_03624_),
    .X(_03626_));
 sg13g2_nor3_1 _09274_ (.A(_03623_),
    .B(_03625_),
    .C(_03626_),
    .Y(_00017_));
 sg13g2_nor2_1 _09275_ (.A(\uart0.rxdiv[3] ),
    .B(_03626_),
    .Y(_03627_));
 sg13g2_and2_1 _09276_ (.A(\uart0.rxdiv[3] ),
    .B(_03626_),
    .X(_03628_));
 sg13g2_nor3_1 _09277_ (.A(_03623_),
    .B(_03627_),
    .C(_03628_),
    .Y(_00018_));
 sg13g2_nand2_1 _09278_ (.Y(_03629_),
    .A(\uart0.rxdiv[4] ),
    .B(_03628_));
 sg13g2_a21oi_1 _09279_ (.A1(\uart0.rxdiv[4] ),
    .A2(_03628_),
    .Y(_03630_),
    .B1(_03623_));
 sg13g2_o21ai_1 _09280_ (.B1(_03630_),
    .Y(_03631_),
    .A1(\uart0.rxdiv[4] ),
    .A2(_03628_));
 sg13g2_inv_1 _09281_ (.Y(_00019_),
    .A(_03631_));
 sg13g2_xor2_1 _09282_ (.B(_03629_),
    .A(\uart0.rxdiv[5] ),
    .X(_03632_));
 sg13g2_nor2_1 _09283_ (.A(_03623_),
    .B(_03632_),
    .Y(_00020_));
 sg13g2_nor2b_1 _09284_ (.A(net3927),
    .B_N(\jtag0.tapst[2] ),
    .Y(_03633_));
 sg13g2_nand2_2 _09285_ (.Y(_03634_),
    .A(net3927),
    .B(_01699_));
 sg13g2_nor2_1 _09286_ (.A(_02550_),
    .B(_03634_),
    .Y(_03635_));
 sg13g2_a21oi_1 _09287_ (.A1(_01748_),
    .A2(_03635_),
    .Y(_03636_),
    .B1(_03633_));
 sg13g2_nor3_1 _09288_ (.A(\jtag0.tapst[3] ),
    .B(\jtag0.tapst[2] ),
    .C(_03634_),
    .Y(_03637_));
 sg13g2_nor2_1 _09289_ (.A(_03378_),
    .B(_03634_),
    .Y(_03638_));
 sg13g2_nor3_1 _09290_ (.A(_01749_),
    .B(_03378_),
    .C(_03634_),
    .Y(_03639_));
 sg13g2_o21ai_1 _09291_ (.B1(_02551_),
    .Y(_03640_),
    .A1(net3926),
    .A2(_03380_));
 sg13g2_nor2_1 _09292_ (.A(_01748_),
    .B(_02585_),
    .Y(_03641_));
 sg13g2_a22oi_1 _09293_ (.Y(_03642_),
    .B1(_02586_),
    .B2(_01748_),
    .A2(_01751_),
    .A1(_00124_));
 sg13g2_a221oi_1 _09294_ (.B2(_03641_),
    .C1(_03639_),
    .B1(_03640_),
    .A1(\jtag0.stms ),
    .Y(_03643_),
    .A2(_03637_));
 sg13g2_nand3_1 _09295_ (.B(_03642_),
    .C(_03643_),
    .A(_03636_),
    .Y(_01535_));
 sg13g2_nor3_1 _09296_ (.A(\jtag0.stms ),
    .B(_01750_),
    .C(_03634_),
    .Y(_03644_));
 sg13g2_a221oi_1 _09297_ (.B2(_00124_),
    .C1(_03644_),
    .B1(_03637_),
    .A1(\jtag0.tapst[1] ),
    .Y(_03645_),
    .A2(_03633_));
 sg13g2_nor2_1 _09298_ (.A(_03378_),
    .B(_03380_),
    .Y(_03646_));
 sg13g2_o21ai_1 _09299_ (.B1(_01749_),
    .Y(_03647_),
    .A1(_03635_),
    .A2(_03646_));
 sg13g2_nor2_1 _09300_ (.A(_02550_),
    .B(_03380_),
    .Y(_03648_));
 sg13g2_o21ai_1 _09301_ (.B1(\jtag0.stms ),
    .Y(_03649_),
    .A1(_03638_),
    .A2(_03648_));
 sg13g2_nand4_1 _09302_ (.B(_03645_),
    .C(_03647_),
    .A(_03642_),
    .Y(_01536_),
    .D(_03649_));
 sg13g2_o21ai_1 _09303_ (.B1(\jtag0.tapst[1] ),
    .Y(_03650_),
    .A1(_02585_),
    .A2(_03633_));
 sg13g2_a22oi_1 _09304_ (.Y(_03651_),
    .B1(\jtag0.stms ),
    .B2(_01751_),
    .A2(net3926),
    .A1(_01699_));
 sg13g2_o21ai_1 _09305_ (.B1(_03651_),
    .Y(_01537_),
    .A1(_00124_),
    .A2(_03650_));
 sg13g2_nand2b_1 _09306_ (.Y(_03652_),
    .B(_01752_),
    .A_N(_03378_));
 sg13g2_a221oi_1 _09307_ (.B2(_00124_),
    .C1(_01751_),
    .B1(_03640_),
    .A1(\jtag0.stms ),
    .Y(_03653_),
    .A2(_03637_));
 sg13g2_nand3b_1 _09308_ (.B(_03652_),
    .C(_03653_),
    .Y(_01538_),
    .A_N(_03644_));
 sg13g2_nor2_1 _09309_ (.A(\cpu.IR[5] ),
    .B(net3393),
    .Y(_03654_));
 sg13g2_nand2b_2 _09310_ (.Y(_03655_),
    .B(net3438),
    .A_N(\cpu.IR[5] ));
 sg13g2_nand2_1 _09311_ (.Y(_03656_),
    .A(\cpu.PCci[31] ),
    .B(net3363));
 sg13g2_o21ai_1 _09312_ (.B1(_03656_),
    .Y(_03657_),
    .A1(_02382_),
    .A2(net3436));
 sg13g2_nand2_1 _09313_ (.Y(_03658_),
    .A(net3367),
    .B(_02647_));
 sg13g2_or3_1 _09314_ (.A(net3451),
    .B(_01762_),
    .C(net3423),
    .X(_03659_));
 sg13g2_o21ai_1 _09315_ (.B1(net3644),
    .Y(_03660_),
    .A1(net3438),
    .A2(net3385));
 sg13g2_nand2_2 _09316_ (.Y(_03661_),
    .A(_03658_),
    .B(_03660_));
 sg13g2_xnor2_1 _09317_ (.Y(_03662_),
    .A(net3335),
    .B(_03661_));
 sg13g2_nand2_1 _09318_ (.Y(_03663_),
    .A(_03657_),
    .B(_03662_));
 sg13g2_xnor2_1 _09319_ (.Y(_03664_),
    .A(_03657_),
    .B(_03662_));
 sg13g2_a22oi_1 _09320_ (.Y(_03665_),
    .B1(net3363),
    .B2(\cpu.PCci[30] ),
    .A2(net3392),
    .A1(_01791_));
 sg13g2_inv_1 _09321_ (.Y(_03666_),
    .A(_03665_));
 sg13g2_and2_1 _09322_ (.A(net3644),
    .B(net3385),
    .X(_03667_));
 sg13g2_nand2_1 _09323_ (.Y(_03668_),
    .A(net3644),
    .B(net3385));
 sg13g2_a22oi_1 _09324_ (.Y(_03669_),
    .B1(net3366),
    .B2(_02743_),
    .A2(net3436),
    .A1(\cpu.Bimm[10] ));
 sg13g2_nand2_2 _09325_ (.Y(_03670_),
    .A(net3360),
    .B(_03669_));
 sg13g2_xnor2_1 _09326_ (.Y(_03671_),
    .A(net3332),
    .B(_03670_));
 sg13g2_nor2_1 _09327_ (.A(_03665_),
    .B(_03671_),
    .Y(_03672_));
 sg13g2_xnor2_1 _09328_ (.Y(_03673_),
    .A(_03666_),
    .B(_03671_));
 sg13g2_nor2_2 _09329_ (.A(_00564_),
    .B(_03655_),
    .Y(_03674_));
 sg13g2_a21oi_2 _09330_ (.B1(_03674_),
    .Y(_03675_),
    .A2(net3394),
    .A1(_01905_));
 sg13g2_a21o_1 _09331_ (.A2(net3394),
    .A1(_01905_),
    .B1(_03674_),
    .X(_03676_));
 sg13g2_nand4_1 _09332_ (.B(_03006_),
    .C(_03008_),
    .A(_02444_),
    .Y(_03677_),
    .D(_03013_));
 sg13g2_a22oi_1 _09333_ (.Y(_03678_),
    .B1(_02473_),
    .B2(\cpu.IR[23] ),
    .A2(net3451),
    .A1(\cpu.Bimm[3] ));
 sg13g2_and2_1 _09334_ (.A(_03677_),
    .B(_03678_),
    .X(_03679_));
 sg13g2_nand2_1 _09335_ (.Y(_03680_),
    .A(_03677_),
    .B(_03678_));
 sg13g2_nand3_1 _09336_ (.B(_03677_),
    .C(_03678_),
    .A(net3336),
    .Y(_03681_));
 sg13g2_a21o_1 _09337_ (.A2(_03678_),
    .A1(_03677_),
    .B1(net3336),
    .X(_03682_));
 sg13g2_a21oi_1 _09338_ (.A1(_03681_),
    .A2(_03682_),
    .Y(_03683_),
    .B1(_03676_));
 sg13g2_a21o_1 _09339_ (.A2(_03682_),
    .A1(_03681_),
    .B1(_03676_),
    .X(_03684_));
 sg13g2_nand2_1 _09340_ (.Y(_03685_),
    .A(_01725_),
    .B(net3365));
 sg13g2_a22oi_1 _09341_ (.Y(_03686_),
    .B1(net3365),
    .B2(_01725_),
    .A2(net3393),
    .A1(_01926_));
 sg13g2_o21ai_1 _09342_ (.B1(_03685_),
    .Y(_03687_),
    .A1(_01927_),
    .A2(net3438));
 sg13g2_nand4_1 _09343_ (.B(_03093_),
    .C(_03095_),
    .A(net3368),
    .Y(_03688_),
    .D(_03100_));
 sg13g2_a22oi_1 _09344_ (.Y(_03689_),
    .B1(_02473_),
    .B2(\cpu.IR[22] ),
    .A2(net3451),
    .A1(\cpu.Bimm[2] ));
 sg13g2_and2_1 _09345_ (.A(_03688_),
    .B(_03689_),
    .X(_03690_));
 sg13g2_nand2_1 _09346_ (.Y(_03691_),
    .A(_03688_),
    .B(_03689_));
 sg13g2_and3_1 _09347_ (.X(_03692_),
    .A(net3336),
    .B(_03688_),
    .C(_03689_));
 sg13g2_a21oi_1 _09348_ (.A1(_03688_),
    .A2(_03689_),
    .Y(_03693_),
    .B1(net3335));
 sg13g2_nor3_1 _09349_ (.A(_03686_),
    .B(_03692_),
    .C(_03693_),
    .Y(_03694_));
 sg13g2_or3_1 _09350_ (.A(_03686_),
    .B(_03692_),
    .C(_03693_),
    .X(_03695_));
 sg13g2_nand3_1 _09351_ (.B(_03681_),
    .C(_03682_),
    .A(_03676_),
    .Y(_03696_));
 sg13g2_o21ai_1 _09352_ (.B1(_02479_),
    .Y(_03697_),
    .A1(_02480_),
    .A2(_02503_));
 sg13g2_o21ai_1 _09353_ (.B1(_03686_),
    .Y(_03698_),
    .A1(_03692_),
    .A2(_03693_));
 sg13g2_and2_1 _09354_ (.A(_03695_),
    .B(_03698_),
    .X(_03699_));
 sg13g2_nand2_1 _09355_ (.Y(_03700_),
    .A(_03684_),
    .B(_03696_));
 sg13g2_and4_1 _09356_ (.A(_03684_),
    .B(_03695_),
    .C(_03696_),
    .D(_03698_),
    .X(_03701_));
 sg13g2_a21oi_1 _09357_ (.A1(_03695_),
    .A2(_03696_),
    .Y(_03702_),
    .B1(_03683_));
 sg13g2_a21o_1 _09358_ (.A2(_03701_),
    .A1(_03697_),
    .B1(_03702_),
    .X(_03703_));
 sg13g2_a21oi_2 _09359_ (.B1(_03702_),
    .Y(_03704_),
    .A2(_03701_),
    .A1(_03697_));
 sg13g2_and2_1 _09360_ (.A(\cpu.PCci[7] ),
    .B(net3365),
    .X(_03705_));
 sg13g2_a21oi_1 _09361_ (.A1(_01855_),
    .A2(net3394),
    .Y(_03706_),
    .B1(_03705_));
 sg13g2_a21o_2 _09362_ (.A2(net3394),
    .A1(_01855_),
    .B1(_03705_),
    .X(_03707_));
 sg13g2_nand3_1 _09363_ (.B(_02656_),
    .C(_02662_),
    .A(net3368),
    .Y(_03708_));
 sg13g2_nand2_1 _09364_ (.Y(_03709_),
    .A(\cpu.Bimm[7] ),
    .B(_03659_));
 sg13g2_nand2_1 _09365_ (.Y(_03710_),
    .A(_03708_),
    .B(_03709_));
 sg13g2_and3_1 _09366_ (.X(_03711_),
    .A(net3334),
    .B(_03708_),
    .C(_03709_));
 sg13g2_a21oi_1 _09367_ (.A1(_03708_),
    .A2(_03709_),
    .Y(_03712_),
    .B1(net3334));
 sg13g2_o21ai_1 _09368_ (.B1(_03707_),
    .Y(_03713_),
    .A1(_03711_),
    .A2(_03712_));
 sg13g2_nor3_1 _09369_ (.A(_03707_),
    .B(_03711_),
    .C(_03712_),
    .Y(_03714_));
 sg13g2_or3_1 _09370_ (.A(_03707_),
    .B(_03711_),
    .C(_03712_),
    .X(_03715_));
 sg13g2_nand2_1 _09371_ (.Y(_03716_),
    .A(_03713_),
    .B(_03715_));
 sg13g2_nor2_1 _09372_ (.A(_00566_),
    .B(_03655_),
    .Y(_03717_));
 sg13g2_a21o_2 _09373_ (.A2(net3394),
    .A1(_01994_),
    .B1(_03717_),
    .X(_03718_));
 sg13g2_nand3_1 _09374_ (.B(_02752_),
    .C(_02758_),
    .A(net3368),
    .Y(_03719_));
 sg13g2_nand2_1 _09375_ (.Y(_03720_),
    .A(\cpu.Bimm[6] ),
    .B(net3385));
 sg13g2_nand2_1 _09376_ (.Y(_03721_),
    .A(_03719_),
    .B(_03720_));
 sg13g2_and3_1 _09377_ (.X(_03722_),
    .A(net3334),
    .B(_03719_),
    .C(_03720_));
 sg13g2_a21oi_1 _09378_ (.A1(_03719_),
    .A2(_03720_),
    .Y(_03723_),
    .B1(net3333));
 sg13g2_o21ai_1 _09379_ (.B1(_03718_),
    .Y(_03724_),
    .A1(_03722_),
    .A2(_03723_));
 sg13g2_or3_1 _09380_ (.A(_03718_),
    .B(_03722_),
    .C(_03723_),
    .X(_03725_));
 sg13g2_nand2_2 _09381_ (.Y(_03726_),
    .A(_03724_),
    .B(_03725_));
 sg13g2_and4_1 _09382_ (.A(_03713_),
    .B(_03715_),
    .C(_03724_),
    .D(_03725_),
    .X(_03727_));
 sg13g2_and2_1 _09383_ (.A(\cpu.PCci[5] ),
    .B(net3365),
    .X(_03728_));
 sg13g2_a21o_2 _09384_ (.A2(net3395),
    .A1(_01871_),
    .B1(_03728_),
    .X(_03729_));
 sg13g2_nand3_1 _09385_ (.B(_02835_),
    .C(_02841_),
    .A(net3368),
    .Y(_03730_));
 sg13g2_nand2_1 _09386_ (.Y(_03731_),
    .A(\cpu.Bimm[5] ),
    .B(net3385));
 sg13g2_nand2_1 _09387_ (.Y(_03732_),
    .A(_03730_),
    .B(_03731_));
 sg13g2_and3_1 _09388_ (.X(_03733_),
    .A(net3333),
    .B(_03730_),
    .C(_03731_));
 sg13g2_a21oi_1 _09389_ (.A1(_03730_),
    .A2(_03731_),
    .Y(_03734_),
    .B1(net3333));
 sg13g2_nor3_1 _09390_ (.A(_03729_),
    .B(_03733_),
    .C(_03734_),
    .Y(_03735_));
 sg13g2_o21ai_1 _09391_ (.B1(_03729_),
    .Y(_03736_),
    .A1(_03733_),
    .A2(_03734_));
 sg13g2_nand2b_1 _09392_ (.Y(_03737_),
    .B(_03736_),
    .A_N(_03735_));
 sg13g2_nor2_1 _09393_ (.A(_00565_),
    .B(_03655_),
    .Y(_03738_));
 sg13g2_a21oi_2 _09394_ (.B1(_03738_),
    .Y(_03739_),
    .A2(net3395),
    .A1(_01887_));
 sg13g2_a21o_1 _09395_ (.A2(net3395),
    .A1(_01887_),
    .B1(_03738_),
    .X(_03740_));
 sg13g2_and3_1 _09396_ (.X(_03741_),
    .A(net3368),
    .B(_02920_),
    .C(_02926_));
 sg13g2_nand2_1 _09397_ (.Y(_03742_),
    .A(\cpu.Bimm[4] ),
    .B(net3451));
 sg13g2_nand2_1 _09398_ (.Y(_03743_),
    .A(\cpu.IR[24] ),
    .B(_02473_));
 sg13g2_and2_1 _09399_ (.A(_03742_),
    .B(_03743_),
    .X(_03744_));
 sg13g2_nand2_1 _09400_ (.Y(_03745_),
    .A(_03742_),
    .B(_03743_));
 sg13g2_nor2_1 _09401_ (.A(_03741_),
    .B(_03745_),
    .Y(_03746_));
 sg13g2_nand2b_1 _09402_ (.Y(_03747_),
    .B(_03744_),
    .A_N(_03741_));
 sg13g2_o21ai_1 _09403_ (.B1(net3333),
    .Y(_03748_),
    .A1(_03741_),
    .A2(_03745_));
 sg13g2_nand3b_1 _09404_ (.B(_03744_),
    .C(net3336),
    .Y(_03749_),
    .A_N(_03741_));
 sg13g2_nand2_1 _09405_ (.Y(_03750_),
    .A(_03748_),
    .B(_03749_));
 sg13g2_nand3_1 _09406_ (.B(_03748_),
    .C(_03749_),
    .A(_03740_),
    .Y(_03751_));
 sg13g2_xnor2_1 _09407_ (.Y(_03752_),
    .A(_03739_),
    .B(_03750_));
 sg13g2_nor4_1 _09408_ (.A(_03716_),
    .B(_03726_),
    .C(_03737_),
    .D(_03752_),
    .Y(_03753_));
 sg13g2_or4_1 _09409_ (.A(_03716_),
    .B(_03726_),
    .C(_03737_),
    .D(_03752_),
    .X(_03754_));
 sg13g2_and2_1 _09410_ (.A(_03736_),
    .B(_03751_),
    .X(_03755_));
 sg13g2_a21oi_1 _09411_ (.A1(_03736_),
    .A2(_03751_),
    .Y(_03756_),
    .B1(_03735_));
 sg13g2_o21ai_1 _09412_ (.B1(_03713_),
    .Y(_03757_),
    .A1(_03714_),
    .A2(_03724_));
 sg13g2_a21oi_1 _09413_ (.A1(_03727_),
    .A2(_03756_),
    .Y(_03758_),
    .B1(_03757_));
 sg13g2_a221oi_1 _09414_ (.B2(_03727_),
    .C1(_03757_),
    .B1(_03756_),
    .A1(_03703_),
    .Y(_03759_),
    .A2(_03753_));
 sg13g2_o21ai_1 _09415_ (.B1(_03758_),
    .Y(_03760_),
    .A1(_03704_),
    .A2(_03754_));
 sg13g2_and2_1 _09416_ (.A(\cpu.PCci[14] ),
    .B(net3364),
    .X(_03761_));
 sg13g2_a21o_2 _09417_ (.A2(net3392),
    .A1(_01824_),
    .B1(_03761_),
    .X(_03762_));
 sg13g2_a21oi_1 _09418_ (.A1(net3694),
    .A2(net3436),
    .Y(_03763_),
    .B1(net3361));
 sg13g2_o21ai_1 _09419_ (.B1(_03763_),
    .Y(_03764_),
    .A1(net3369),
    .A2(_02776_));
 sg13g2_xnor2_1 _09420_ (.Y(_03765_),
    .A(net3332),
    .B(_03764_));
 sg13g2_nor2b_1 _09421_ (.A(_03765_),
    .B_N(_03762_),
    .Y(_03766_));
 sg13g2_nand2b_1 _09422_ (.Y(_03767_),
    .B(_03762_),
    .A_N(_03765_));
 sg13g2_xor2_1 _09423_ (.B(_03765_),
    .A(_03762_),
    .X(_03768_));
 sg13g2_a22oi_1 _09424_ (.Y(_03769_),
    .B1(net3364),
    .B2(\cpu.PCci[15] ),
    .A2(net3392),
    .A1(_01807_));
 sg13g2_a21oi_1 _09425_ (.A1(net3680),
    .A2(net3437),
    .Y(_03770_),
    .B1(net3361));
 sg13g2_o21ai_1 _09426_ (.B1(_03770_),
    .Y(_03771_),
    .A1(net3369),
    .A2(_02680_));
 sg13g2_inv_1 _09427_ (.Y(_03772_),
    .A(_03771_));
 sg13g2_xnor2_1 _09428_ (.Y(_03773_),
    .A(net3332),
    .B(_03771_));
 sg13g2_nor2_1 _09429_ (.A(_03769_),
    .B(_03773_),
    .Y(_03774_));
 sg13g2_nand2_1 _09430_ (.Y(_03775_),
    .A(_03769_),
    .B(_03773_));
 sg13g2_xnor2_1 _09431_ (.Y(_03776_),
    .A(_03769_),
    .B(_03773_));
 sg13g2_or2_1 _09432_ (.X(_03777_),
    .B(_03776_),
    .A(_03768_));
 sg13g2_a22oi_1 _09433_ (.Y(_03778_),
    .B1(net3364),
    .B2(\cpu.PCci[13] ),
    .A2(net3392),
    .A1(_02097_));
 sg13g2_a21oi_1 _09434_ (.A1(net3697),
    .A2(net3436),
    .Y(_03779_),
    .B1(net3361));
 sg13g2_o21ai_1 _09435_ (.B1(_03779_),
    .Y(_03780_),
    .A1(net3369),
    .A2(_02859_));
 sg13g2_inv_1 _09436_ (.Y(_03781_),
    .A(_03780_));
 sg13g2_xnor2_1 _09437_ (.Y(_03782_),
    .A(net3332),
    .B(_03780_));
 sg13g2_nand2_1 _09438_ (.Y(_03783_),
    .A(_03778_),
    .B(_03782_));
 sg13g2_nor2_1 _09439_ (.A(_03778_),
    .B(_03782_),
    .Y(_03784_));
 sg13g2_xnor2_1 _09440_ (.Y(_03785_),
    .A(_03778_),
    .B(_03782_));
 sg13g2_a22oi_1 _09441_ (.Y(_03786_),
    .B1(net3364),
    .B2(_01728_),
    .A2(net3392),
    .A1(_02078_));
 sg13g2_a21oi_1 _09442_ (.A1(\cpu.IR[12] ),
    .A2(net3436),
    .Y(_03787_),
    .B1(net3361));
 sg13g2_o21ai_1 _09443_ (.B1(_03787_),
    .Y(_03788_),
    .A1(net3369),
    .A2(_02945_));
 sg13g2_inv_1 _09444_ (.Y(_03789_),
    .A(_03788_));
 sg13g2_xnor2_1 _09445_ (.Y(_03790_),
    .A(net3332),
    .B(_03788_));
 sg13g2_nor2_1 _09446_ (.A(_03786_),
    .B(_03790_),
    .Y(_03791_));
 sg13g2_xnor2_1 _09447_ (.Y(_03792_),
    .A(_03786_),
    .B(_03790_));
 sg13g2_nor4_2 _09448_ (.A(_03768_),
    .B(_03776_),
    .C(_03785_),
    .Y(_03793_),
    .D(_03792_));
 sg13g2_a22oi_1 _09449_ (.Y(_03794_),
    .B1(net3365),
    .B2(_01727_),
    .A2(net3393),
    .A1(_02053_));
 sg13g2_nand2_1 _09450_ (.Y(_03795_),
    .A(\cpu.Bimm[10] ),
    .B(net3385));
 sg13g2_o21ai_1 _09451_ (.B1(_03795_),
    .Y(_03796_),
    .A1(net3369),
    .A2(_03118_));
 sg13g2_inv_1 _09452_ (.Y(_03797_),
    .A(_03796_));
 sg13g2_xnor2_1 _09453_ (.Y(_03798_),
    .A(net3333),
    .B(_03796_));
 sg13g2_nor2_1 _09454_ (.A(_03794_),
    .B(_03798_),
    .Y(_03799_));
 sg13g2_xor2_1 _09455_ (.B(_03798_),
    .A(_03794_),
    .X(_03800_));
 sg13g2_and2_1 _09456_ (.A(_01839_),
    .B(net3394),
    .X(_03801_));
 sg13g2_a21oi_2 _09457_ (.B1(_03801_),
    .Y(_03802_),
    .A2(_03654_),
    .A1(\cpu.PCci[11] ));
 sg13g2_a21o_2 _09458_ (.A2(net3365),
    .A1(\cpu.PCci[11] ),
    .B1(_03801_),
    .X(_03803_));
 sg13g2_o21ai_1 _09459_ (.B1(net3360),
    .Y(_03804_),
    .A1(net3370),
    .A2(_03031_));
 sg13g2_xnor2_1 _09460_ (.Y(_03805_),
    .A(net3335),
    .B(_03804_));
 sg13g2_nand2b_1 _09461_ (.Y(_03806_),
    .B(_03802_),
    .A_N(_03805_));
 sg13g2_and2_1 _09462_ (.A(_03803_),
    .B(_03805_),
    .X(_03807_));
 sg13g2_xnor2_1 _09463_ (.Y(_03808_),
    .A(_03802_),
    .B(_03805_));
 sg13g2_and2_1 _09464_ (.A(_03800_),
    .B(_03808_),
    .X(_03809_));
 sg13g2_nand2_1 _09465_ (.Y(_03810_),
    .A(_03800_),
    .B(_03808_));
 sg13g2_nand2_1 _09466_ (.Y(_03811_),
    .A(_02014_),
    .B(net3393));
 sg13g2_o21ai_1 _09467_ (.B1(_03811_),
    .Y(_03812_),
    .A1(_00567_),
    .A2(_03655_));
 sg13g2_nand2_1 _09468_ (.Y(_03813_),
    .A(\cpu.Bimm[8] ),
    .B(net3385));
 sg13g2_o21ai_1 _09469_ (.B1(_03813_),
    .Y(_03814_),
    .A1(net3370),
    .A2(_03265_));
 sg13g2_xnor2_1 _09470_ (.Y(_03815_),
    .A(net3333),
    .B(_03814_));
 sg13g2_nor2b_1 _09471_ (.A(_03815_),
    .B_N(_03812_),
    .Y(_03816_));
 sg13g2_xnor2_1 _09472_ (.Y(_03817_),
    .A(_03812_),
    .B(_03815_));
 sg13g2_inv_1 _09473_ (.Y(_03818_),
    .A(_03817_));
 sg13g2_a22oi_1 _09474_ (.Y(_03819_),
    .B1(net3365),
    .B2(\cpu.PCci[9] ),
    .A2(net3393),
    .A1(_02033_));
 sg13g2_nand4_1 _09475_ (.B(_03183_),
    .C(_03185_),
    .A(net3368),
    .Y(_03820_),
    .D(_03190_));
 sg13g2_nand2_1 _09476_ (.Y(_03821_),
    .A(\cpu.Bimm[9] ),
    .B(net3385));
 sg13g2_and2_1 _09477_ (.A(_03820_),
    .B(_03821_),
    .X(_03822_));
 sg13g2_xnor2_1 _09478_ (.Y(_03823_),
    .A(net3335),
    .B(_03822_));
 sg13g2_nand2_1 _09479_ (.Y(_03824_),
    .A(_03819_),
    .B(_03823_));
 sg13g2_nor2_1 _09480_ (.A(_03819_),
    .B(_03823_),
    .Y(_03825_));
 sg13g2_xor2_1 _09481_ (.B(_03823_),
    .A(_03819_),
    .X(_03826_));
 sg13g2_and4_1 _09482_ (.A(_03793_),
    .B(_03809_),
    .C(_03817_),
    .D(_03826_),
    .X(_03827_));
 sg13g2_a21oi_2 _09483_ (.B1(_03807_),
    .Y(_03828_),
    .A2(_03806_),
    .A1(_03799_));
 sg13g2_nor2_1 _09484_ (.A(_03816_),
    .B(_03825_),
    .Y(_03829_));
 sg13g2_o21ai_1 _09485_ (.B1(_03824_),
    .Y(_03830_),
    .A1(_03816_),
    .A2(_03825_));
 sg13g2_o21ai_1 _09486_ (.B1(_03828_),
    .Y(_03831_),
    .A1(_03810_),
    .A2(_03830_));
 sg13g2_a21oi_1 _09487_ (.A1(_03766_),
    .A2(_03775_),
    .Y(_03832_),
    .B1(_03774_));
 sg13g2_or2_1 _09488_ (.X(_03833_),
    .B(_03791_),
    .A(_03784_));
 sg13g2_a21oi_1 _09489_ (.A1(_03783_),
    .A2(_03791_),
    .Y(_03834_),
    .B1(_03784_));
 sg13g2_o21ai_1 _09490_ (.B1(_03832_),
    .Y(_03835_),
    .A1(_03777_),
    .A2(_03834_));
 sg13g2_a221oi_1 _09491_ (.B2(_03793_),
    .C1(_03835_),
    .B1(_03831_),
    .A1(_03760_),
    .Y(_03836_),
    .A2(_03827_));
 sg13g2_a22oi_1 _09492_ (.Y(_03837_),
    .B1(net3363),
    .B2(\cpu.PCci[19] ),
    .A2(net3392),
    .A1(_02242_));
 sg13g2_a21oi_1 _09493_ (.A1(\cpu.IR[19] ),
    .A2(net3436),
    .Y(_03838_),
    .B1(net3361));
 sg13g2_o21ai_1 _09494_ (.B1(_03838_),
    .Y(_03839_),
    .A1(net3369),
    .A2(_03052_));
 sg13g2_inv_1 _09495_ (.Y(_03840_),
    .A(_03839_));
 sg13g2_xnor2_1 _09496_ (.Y(_03841_),
    .A(net3331),
    .B(_03839_));
 sg13g2_nor2_1 _09497_ (.A(_03837_),
    .B(_03841_),
    .Y(_03842_));
 sg13g2_nand2_1 _09498_ (.Y(_03843_),
    .A(_03837_),
    .B(_03841_));
 sg13g2_xnor2_1 _09499_ (.Y(_03844_),
    .A(_03837_),
    .B(_03841_));
 sg13g2_inv_1 _09500_ (.Y(_03845_),
    .A(_03844_));
 sg13g2_and2_1 _09501_ (.A(\cpu.PCci[18] ),
    .B(net3362),
    .X(_03846_));
 sg13g2_a21o_2 _09502_ (.A2(net3391),
    .A1(_02205_),
    .B1(_03846_),
    .X(_03847_));
 sg13g2_a21oi_1 _09503_ (.A1(\cpu.IR[18] ),
    .A2(net3435),
    .Y(_03848_),
    .B1(net3361));
 sg13g2_o21ai_1 _09504_ (.B1(_03848_),
    .Y(_03849_),
    .A1(net3369),
    .A2(_03140_));
 sg13g2_xnor2_1 _09505_ (.Y(_03850_),
    .A(net3332),
    .B(_03849_));
 sg13g2_nor2b_1 _09506_ (.A(_03850_),
    .B_N(_03847_),
    .Y(_03851_));
 sg13g2_xor2_1 _09507_ (.B(_03850_),
    .A(_03847_),
    .X(_03852_));
 sg13g2_or2_1 _09508_ (.X(_03853_),
    .B(_03852_),
    .A(_03844_));
 sg13g2_a22oi_1 _09509_ (.Y(_03854_),
    .B1(net3364),
    .B2(\cpu.PCci[17] ),
    .A2(net3391),
    .A1(_02222_));
 sg13g2_a21oi_1 _09510_ (.A1(net3655),
    .A2(net3435),
    .Y(_03855_),
    .B1(net3361));
 sg13g2_o21ai_1 _09511_ (.B1(_03855_),
    .Y(_03856_),
    .A1(net3369),
    .A2(_03214_));
 sg13g2_inv_1 _09512_ (.Y(_03857_),
    .A(_03856_));
 sg13g2_xnor2_1 _09513_ (.Y(_03858_),
    .A(net3332),
    .B(_03856_));
 sg13g2_nand2_1 _09514_ (.Y(_03859_),
    .A(_03854_),
    .B(_03858_));
 sg13g2_nor2_1 _09515_ (.A(_03854_),
    .B(_03858_),
    .Y(_03860_));
 sg13g2_xnor2_1 _09516_ (.Y(_03861_),
    .A(_03854_),
    .B(_03858_));
 sg13g2_nor2_1 _09517_ (.A(_03853_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_a22oi_1 _09518_ (.Y(_03863_),
    .B1(net3362),
    .B2(\cpu.PCci[21] ),
    .A2(net3390),
    .A1(_02171_));
 sg13g2_inv_1 _09519_ (.Y(_03864_),
    .A(_03863_));
 sg13g2_a22oi_1 _09520_ (.Y(_03865_),
    .B1(net3366),
    .B2(_02879_),
    .A2(net3435),
    .A1(\cpu.IR[21] ));
 sg13g2_nand2_2 _09521_ (.Y(_03866_),
    .A(net3359),
    .B(_03865_));
 sg13g2_xnor2_1 _09522_ (.Y(_03867_),
    .A(net3331),
    .B(_03866_));
 sg13g2_nand2b_1 _09523_ (.Y(_03868_),
    .B(_03864_),
    .A_N(_03867_));
 sg13g2_and2_1 _09524_ (.A(_03863_),
    .B(_03867_),
    .X(_03869_));
 sg13g2_xnor2_1 _09525_ (.Y(_03870_),
    .A(_03863_),
    .B(_03867_));
 sg13g2_a22oi_1 _09526_ (.Y(_03871_),
    .B1(net3362),
    .B2(\cpu.PCci[20] ),
    .A2(net3390),
    .A1(_02185_));
 sg13g2_a22oi_1 _09527_ (.Y(_03872_),
    .B1(net3367),
    .B2(_02965_),
    .A2(net3435),
    .A1(net3647));
 sg13g2_nand2_1 _09528_ (.Y(_03873_),
    .A(net3359),
    .B(_03872_));
 sg13g2_xnor2_1 _09529_ (.Y(_03874_),
    .A(net3331),
    .B(_03873_));
 sg13g2_or2_1 _09530_ (.X(_03875_),
    .B(_03874_),
    .A(_03871_));
 sg13g2_xor2_1 _09531_ (.B(_03874_),
    .A(_03871_),
    .X(_03876_));
 sg13g2_xnor2_1 _09532_ (.Y(_03877_),
    .A(_03871_),
    .B(_03874_));
 sg13g2_and2_1 _09533_ (.A(\cpu.PCci[16] ),
    .B(net3364),
    .X(_03878_));
 sg13g2_a21oi_2 _09534_ (.B1(_03878_),
    .Y(_03879_),
    .A2(net3391),
    .A1(_02118_));
 sg13g2_a21o_1 _09535_ (.A2(net3391),
    .A1(_02118_),
    .B1(_03878_),
    .X(_03880_));
 sg13g2_nand4_1 _09536_ (.B(_03279_),
    .C(_03281_),
    .A(net3368),
    .Y(_03881_),
    .D(_03286_));
 sg13g2_a21oi_1 _09537_ (.A1(net3661),
    .A2(net3435),
    .Y(_03882_),
    .B1(net3361));
 sg13g2_nand2_1 _09538_ (.Y(_03883_),
    .A(_03881_),
    .B(_03882_));
 sg13g2_xnor2_1 _09539_ (.Y(_03884_),
    .A(net3331),
    .B(_03883_));
 sg13g2_nor2_1 _09540_ (.A(_03879_),
    .B(_03884_),
    .Y(_03885_));
 sg13g2_xnor2_1 _09541_ (.Y(_03886_),
    .A(_03880_),
    .B(_03884_));
 sg13g2_xnor2_1 _09542_ (.Y(_03887_),
    .A(_03879_),
    .B(_03884_));
 sg13g2_a22oi_1 _09543_ (.Y(_03888_),
    .B1(net3362),
    .B2(\cpu.PCci[22] ),
    .A2(net3390),
    .A1(_02134_));
 sg13g2_a22oi_1 _09544_ (.Y(_03889_),
    .B1(net3366),
    .B2(_02796_),
    .A2(net3437),
    .A1(\cpu.IR[22] ));
 sg13g2_nand2_2 _09545_ (.Y(_03890_),
    .A(net3359),
    .B(_03889_));
 sg13g2_xnor2_1 _09546_ (.Y(_03891_),
    .A(net3331),
    .B(_03890_));
 sg13g2_nor2_1 _09547_ (.A(_03888_),
    .B(_03891_),
    .Y(_03892_));
 sg13g2_nand2_1 _09548_ (.Y(_03893_),
    .A(_03888_),
    .B(_03891_));
 sg13g2_xnor2_1 _09549_ (.Y(_03894_),
    .A(_03888_),
    .B(_03891_));
 sg13g2_and2_1 _09550_ (.A(\cpu.PCci[23] ),
    .B(net3362),
    .X(_03895_));
 sg13g2_a21o_2 _09551_ (.A2(net3390),
    .A1(_02152_),
    .B1(_03895_),
    .X(_03896_));
 sg13g2_a22oi_1 _09552_ (.Y(_03897_),
    .B1(net3366),
    .B2(_02701_),
    .A2(net3435),
    .A1(\cpu.IR[23] ));
 sg13g2_nand2_2 _09553_ (.Y(_03898_),
    .A(net3359),
    .B(_03897_));
 sg13g2_xnor2_1 _09554_ (.Y(_03899_),
    .A(net3331),
    .B(_03898_));
 sg13g2_nor2b_1 _09555_ (.A(_03899_),
    .B_N(_03896_),
    .Y(_03900_));
 sg13g2_nand2b_1 _09556_ (.Y(_03901_),
    .B(_03899_),
    .A_N(_03896_));
 sg13g2_xor2_1 _09557_ (.B(_03899_),
    .A(_03896_),
    .X(_03902_));
 sg13g2_nor2_1 _09558_ (.A(_03894_),
    .B(_03902_),
    .Y(_03903_));
 sg13g2_nor4_1 _09559_ (.A(_03870_),
    .B(_03877_),
    .C(_03894_),
    .D(_03902_),
    .Y(_03904_));
 sg13g2_nand3_1 _09560_ (.B(_03886_),
    .C(_03904_),
    .A(_03862_),
    .Y(_03905_));
 sg13g2_a21o_1 _09561_ (.A2(_03901_),
    .A1(_03892_),
    .B1(_03900_),
    .X(_03906_));
 sg13g2_a21o_1 _09562_ (.A2(_03875_),
    .A1(_03868_),
    .B1(_03869_),
    .X(_03907_));
 sg13g2_a21oi_1 _09563_ (.A1(_03868_),
    .A2(_03875_),
    .Y(_03908_),
    .B1(_03869_));
 sg13g2_nor2_1 _09564_ (.A(_03860_),
    .B(_03885_),
    .Y(_03909_));
 sg13g2_o21ai_1 _09565_ (.B1(_03859_),
    .Y(_03910_),
    .A1(_03860_),
    .A2(_03885_));
 sg13g2_a21oi_1 _09566_ (.A1(_03843_),
    .A2(_03851_),
    .Y(_03911_),
    .B1(_03842_));
 sg13g2_o21ai_1 _09567_ (.B1(_03911_),
    .Y(_03912_),
    .A1(_03853_),
    .A2(_03910_));
 sg13g2_a221oi_1 _09568_ (.B2(_03904_),
    .C1(_03906_),
    .B1(_03912_),
    .A1(_03903_),
    .Y(_03913_),
    .A2(_03908_));
 sg13g2_o21ai_1 _09569_ (.B1(_03913_),
    .Y(_03914_),
    .A1(_03836_),
    .A2(_03905_));
 sg13g2_and2_1 _09570_ (.A(\cpu.PCci[27] ),
    .B(net3363),
    .X(_03915_));
 sg13g2_a21o_2 _09571_ (.A2(net3390),
    .A1(_02268_),
    .B1(_03915_),
    .X(_03916_));
 sg13g2_inv_1 _09572_ (.Y(_03917_),
    .A(_03916_));
 sg13g2_a22oi_1 _09573_ (.Y(_03918_),
    .B1(net3366),
    .B2(_02997_),
    .A2(net3435),
    .A1(\cpu.Bimm[7] ));
 sg13g2_nand2_2 _09574_ (.Y(_03919_),
    .A(net3359),
    .B(_03918_));
 sg13g2_xnor2_1 _09575_ (.Y(_03920_),
    .A(net3331),
    .B(_03919_));
 sg13g2_nand2_1 _09576_ (.Y(_03921_),
    .A(_03917_),
    .B(_03920_));
 sg13g2_xnor2_1 _09577_ (.Y(_03922_),
    .A(_03916_),
    .B(_03920_));
 sg13g2_a22oi_1 _09578_ (.Y(_03923_),
    .B1(net3362),
    .B2(\cpu.PCci[26] ),
    .A2(net3390),
    .A1(_02282_));
 sg13g2_a22oi_1 _09579_ (.Y(_03924_),
    .B1(net3367),
    .B2(_03084_),
    .A2(net3435),
    .A1(\cpu.Bimm[6] ));
 sg13g2_nand2_1 _09580_ (.Y(_03925_),
    .A(net3359),
    .B(_03924_));
 sg13g2_inv_1 _09581_ (.Y(_03926_),
    .A(_03925_));
 sg13g2_xnor2_1 _09582_ (.Y(_03927_),
    .A(net3331),
    .B(_03925_));
 sg13g2_nor2_1 _09583_ (.A(_03923_),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_xor2_1 _09584_ (.B(_03927_),
    .A(_03923_),
    .X(_03929_));
 sg13g2_a22oi_1 _09585_ (.Y(_03930_),
    .B1(net3362),
    .B2(\cpu.PCci[25] ),
    .A2(net3390),
    .A1(_02314_));
 sg13g2_a221oi_1 _09586_ (.B2(_03174_),
    .C1(_03667_),
    .B1(net3366),
    .A1(\cpu.Bimm[5] ),
    .Y(_03931_),
    .A2(net3437));
 sg13g2_xnor2_1 _09587_ (.Y(_03932_),
    .A(net3335),
    .B(_03931_));
 sg13g2_and2_1 _09588_ (.A(_03930_),
    .B(_03932_),
    .X(_03933_));
 sg13g2_nor2_1 _09589_ (.A(_03930_),
    .B(_03932_),
    .Y(_03934_));
 sg13g2_or2_1 _09590_ (.X(_03935_),
    .B(_03934_),
    .A(_03933_));
 sg13g2_a22oi_1 _09591_ (.Y(_03936_),
    .B1(net3362),
    .B2(\cpu.PCci[24] ),
    .A2(net3390),
    .A1(_02297_));
 sg13g2_a221oi_1 _09592_ (.B2(_03248_),
    .C1(_03667_),
    .B1(net3367),
    .A1(\cpu.IR[24] ),
    .Y(_03937_),
    .A2(net3438));
 sg13g2_xnor2_1 _09593_ (.Y(_03938_),
    .A(net3335),
    .B(_03937_));
 sg13g2_nor2_1 _09594_ (.A(_03936_),
    .B(_03938_),
    .Y(_03939_));
 sg13g2_xor2_1 _09595_ (.B(_03938_),
    .A(_03936_),
    .X(_03940_));
 sg13g2_nand3_1 _09596_ (.B(_03929_),
    .C(_03940_),
    .A(_03922_),
    .Y(_03941_));
 sg13g2_nor2_1 _09597_ (.A(_03935_),
    .B(_03941_),
    .Y(_03942_));
 sg13g2_nor2_1 _09598_ (.A(_03934_),
    .B(_03939_),
    .Y(_03943_));
 sg13g2_nor2_1 _09599_ (.A(_03933_),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_nand3_1 _09600_ (.B(_03929_),
    .C(_03944_),
    .A(_03922_),
    .Y(_03945_));
 sg13g2_o21ai_1 _09601_ (.B1(_03945_),
    .Y(_03946_),
    .A1(_03917_),
    .A2(_03920_));
 sg13g2_a221oi_1 _09602_ (.B2(_03914_),
    .C1(_03946_),
    .B1(_03942_),
    .A1(_03921_),
    .Y(_03947_),
    .A2(_03928_));
 sg13g2_and2_1 _09603_ (.A(_02358_),
    .B(net3392),
    .X(_03948_));
 sg13g2_a21oi_2 _09604_ (.B1(_03948_),
    .Y(_03949_),
    .A2(net3363),
    .A1(\cpu.PCci[29] ));
 sg13g2_a21o_2 _09605_ (.A2(net3363),
    .A1(\cpu.PCci[29] ),
    .B1(_03948_),
    .X(_03950_));
 sg13g2_a22oi_1 _09606_ (.Y(_03951_),
    .B1(net3366),
    .B2(_02826_),
    .A2(net3436),
    .A1(\cpu.Bimm[9] ));
 sg13g2_nand2_2 _09607_ (.Y(_03952_),
    .A(net3360),
    .B(_03951_));
 sg13g2_xnor2_1 _09608_ (.Y(_03953_),
    .A(net3333),
    .B(_03952_));
 sg13g2_inv_1 _09609_ (.Y(_03954_),
    .A(_03953_));
 sg13g2_xnor2_1 _09610_ (.Y(_03955_),
    .A(_03950_),
    .B(_03953_));
 sg13g2_and2_1 _09611_ (.A(\cpu.PCci[28] ),
    .B(net3363),
    .X(_03956_));
 sg13g2_a21o_2 _09612_ (.A2(net3392),
    .A1(_02339_),
    .B1(_03956_),
    .X(_03957_));
 sg13g2_a22oi_1 _09613_ (.Y(_03958_),
    .B1(net3366),
    .B2(_02911_),
    .A2(net3436),
    .A1(\cpu.Bimm[8] ));
 sg13g2_nand2_2 _09614_ (.Y(_03959_),
    .A(net3360),
    .B(_03958_));
 sg13g2_xnor2_1 _09615_ (.Y(_03960_),
    .A(net3332),
    .B(_03959_));
 sg13g2_nand2b_1 _09616_ (.Y(_03961_),
    .B(_03957_),
    .A_N(_03960_));
 sg13g2_xor2_1 _09617_ (.B(_03960_),
    .A(_03957_),
    .X(_03962_));
 sg13g2_inv_1 _09618_ (.Y(_03963_),
    .A(_03962_));
 sg13g2_nand2_1 _09619_ (.Y(_03964_),
    .A(_03955_),
    .B(_03963_));
 sg13g2_a21oi_1 _09620_ (.A1(_03949_),
    .A2(_03953_),
    .Y(_03965_),
    .B1(_03961_));
 sg13g2_a21oi_1 _09621_ (.A1(_03950_),
    .A2(_03954_),
    .Y(_03966_),
    .B1(_03965_));
 sg13g2_o21ai_1 _09622_ (.B1(_03966_),
    .Y(_03967_),
    .A1(_03947_),
    .A2(_03964_));
 sg13g2_a21oi_2 _09623_ (.B1(_03672_),
    .Y(_03968_),
    .A2(_03967_),
    .A1(_03673_));
 sg13g2_o21ai_1 _09624_ (.B1(_03663_),
    .Y(_03969_),
    .A1(_03664_),
    .A2(_03968_));
 sg13g2_xnor2_1 _09625_ (.Y(_03970_),
    .A(net3333),
    .B(_03969_));
 sg13g2_nor2_1 _09626_ (.A(net3624),
    .B(_03970_),
    .Y(_03971_));
 sg13g2_xnor2_1 _09627_ (.Y(_03972_),
    .A(_03657_),
    .B(_03661_));
 sg13g2_a21oi_1 _09628_ (.A1(_03658_),
    .A2(_03660_),
    .Y(_03973_),
    .B1(_03657_));
 sg13g2_a21oi_1 _09629_ (.A1(_03970_),
    .A2(_03972_),
    .Y(_03974_),
    .B1(_03973_));
 sg13g2_a21oi_1 _09630_ (.A1(net3624),
    .A2(_03974_),
    .Y(_03975_),
    .B1(_03971_));
 sg13g2_xnor2_1 _09631_ (.Y(_03976_),
    .A(_01697_),
    .B(_03975_));
 sg13g2_nand2b_1 _09632_ (.Y(_03977_),
    .B(_03886_),
    .A_N(_03836_));
 sg13g2_nor4_1 _09633_ (.A(_03836_),
    .B(_03853_),
    .C(_03861_),
    .D(_03887_),
    .Y(_03978_));
 sg13g2_o21ai_1 _09634_ (.B1(_03876_),
    .Y(_03979_),
    .A1(_03912_),
    .A2(_03978_));
 sg13g2_nand2_1 _09635_ (.Y(_03980_),
    .A(_03875_),
    .B(_03979_));
 sg13g2_o21ai_1 _09636_ (.B1(_03907_),
    .Y(_03981_),
    .A1(_03869_),
    .A2(_03979_));
 sg13g2_a21oi_1 _09637_ (.A1(_03893_),
    .A2(_03981_),
    .Y(_03982_),
    .B1(_03892_));
 sg13g2_xnor2_1 _09638_ (.Y(_03983_),
    .A(_03902_),
    .B(_03982_));
 sg13g2_o21ai_1 _09639_ (.B1(_03829_),
    .Y(_03984_),
    .A1(_03759_),
    .A2(_03818_));
 sg13g2_nand3_1 _09640_ (.B(_03824_),
    .C(_03984_),
    .A(_03800_),
    .Y(_03985_));
 sg13g2_nand3_1 _09641_ (.B(_03824_),
    .C(_03984_),
    .A(_03809_),
    .Y(_03986_));
 sg13g2_a21oi_2 _09642_ (.B1(_03792_),
    .Y(_03987_),
    .A2(_03986_),
    .A1(_03828_));
 sg13g2_o21ai_1 _09643_ (.B1(_03783_),
    .Y(_03988_),
    .A1(_03833_),
    .A2(_03987_));
 sg13g2_o21ai_1 _09644_ (.B1(_03767_),
    .Y(_03989_),
    .A1(_03768_),
    .A2(_03988_));
 sg13g2_xor2_1 _09645_ (.B(_03989_),
    .A(_03776_),
    .X(_03990_));
 sg13g2_xor2_1 _09646_ (.B(_03988_),
    .A(_03768_),
    .X(_03991_));
 sg13g2_nand2_1 _09647_ (.Y(_03992_),
    .A(_03914_),
    .B(_03940_));
 sg13g2_a21oi_1 _09648_ (.A1(_03914_),
    .A2(_03940_),
    .Y(_03993_),
    .B1(_03939_));
 sg13g2_a21oi_1 _09649_ (.A1(_03943_),
    .A2(_03992_),
    .Y(_03994_),
    .B1(_03933_));
 sg13g2_xor2_1 _09650_ (.B(_03994_),
    .A(_03929_),
    .X(_03995_));
 sg13g2_o21ai_1 _09651_ (.B1(_03909_),
    .Y(_03996_),
    .A1(_03836_),
    .A2(_03887_));
 sg13g2_nand2_1 _09652_ (.Y(_03997_),
    .A(_03859_),
    .B(_03996_));
 sg13g2_a221oi_1 _09653_ (.B2(_03977_),
    .C1(_03852_),
    .B1(_03909_),
    .A1(_03854_),
    .Y(_03998_),
    .A2(_03858_));
 sg13g2_xnor2_1 _09654_ (.Y(_03999_),
    .A(_03852_),
    .B(_03997_));
 sg13g2_nor2b_1 _09655_ (.A(_03799_),
    .B_N(_03985_),
    .Y(_04000_));
 sg13g2_xnor2_1 _09656_ (.Y(_04001_),
    .A(_03808_),
    .B(_04000_));
 sg13g2_xor2_1 _09657_ (.B(_04000_),
    .A(_03808_),
    .X(_04002_));
 sg13g2_or3_1 _09658_ (.A(_03876_),
    .B(_03912_),
    .C(_03978_),
    .X(_04003_));
 sg13g2_nand2_2 _09659_ (.Y(_04004_),
    .A(_03979_),
    .B(_04003_));
 sg13g2_and3_1 _09660_ (.X(_04005_),
    .A(_03999_),
    .B(_04002_),
    .C(_04004_));
 sg13g2_o21ai_1 _09661_ (.B1(_03845_),
    .Y(_04006_),
    .A1(_03851_),
    .A2(_03998_));
 sg13g2_or3_1 _09662_ (.A(_03845_),
    .B(_03851_),
    .C(_03998_),
    .X(_04007_));
 sg13g2_nand2_2 _09663_ (.Y(_04008_),
    .A(_04006_),
    .B(_04007_));
 sg13g2_xor2_1 _09664_ (.B(_03980_),
    .A(_03870_),
    .X(_04009_));
 sg13g2_a21oi_1 _09665_ (.A1(_03929_),
    .A2(_03994_),
    .Y(_04010_),
    .B1(_03928_));
 sg13g2_xor2_1 _09666_ (.B(_04010_),
    .A(_03922_),
    .X(_04011_));
 sg13g2_xnor2_1 _09667_ (.Y(_04012_),
    .A(_03894_),
    .B(_03981_));
 sg13g2_xnor2_1 _09668_ (.Y(_04013_),
    .A(_03664_),
    .B(_03968_));
 sg13g2_xor2_1 _09669_ (.B(_03967_),
    .A(_03673_),
    .X(_04014_));
 sg13g2_xnor2_1 _09670_ (.Y(_04015_),
    .A(_03947_),
    .B(_03962_));
 sg13g2_o21ai_1 _09671_ (.B1(_03755_),
    .Y(_04016_),
    .A1(_03704_),
    .A2(_03752_));
 sg13g2_nand2b_1 _09672_ (.Y(_04017_),
    .B(_04016_),
    .A_N(_03735_));
 sg13g2_xor2_1 _09673_ (.B(_04017_),
    .A(_03726_),
    .X(_04018_));
 sg13g2_xnor2_1 _09674_ (.Y(_04019_),
    .A(_03759_),
    .B(_03817_));
 sg13g2_o21ai_1 _09675_ (.B1(_03751_),
    .Y(_04020_),
    .A1(_03704_),
    .A2(_03752_));
 sg13g2_xnor2_1 _09676_ (.Y(_04021_),
    .A(_03737_),
    .B(_04020_));
 sg13g2_a21oi_1 _09677_ (.A1(_03697_),
    .A2(_03699_),
    .Y(_04022_),
    .B1(_03694_));
 sg13g2_xor2_1 _09678_ (.B(_04022_),
    .A(_03700_),
    .X(_04023_));
 sg13g2_xnor2_1 _09679_ (.Y(_04024_),
    .A(_03697_),
    .B(_03699_));
 sg13g2_inv_1 _09680_ (.Y(_04025_),
    .A(_04024_));
 sg13g2_nor4_1 _09681_ (.A(net3140),
    .B(net3236),
    .C(_04023_),
    .D(_04025_),
    .Y(_04026_));
 sg13g2_xnor2_1 _09682_ (.Y(_04027_),
    .A(_03704_),
    .B(_03752_));
 sg13g2_nand3b_1 _09683_ (.B(_04026_),
    .C(_04027_),
    .Y(_04028_),
    .A_N(_04021_));
 sg13g2_a21oi_1 _09684_ (.A1(_03760_),
    .A2(_03817_),
    .Y(_04029_),
    .B1(_03816_));
 sg13g2_xor2_1 _09685_ (.B(_04029_),
    .A(_03826_),
    .X(_04030_));
 sg13g2_xnor2_1 _09686_ (.Y(_04031_),
    .A(_03836_),
    .B(_03886_));
 sg13g2_inv_1 _09687_ (.Y(_04032_),
    .A(_04031_));
 sg13g2_nor4_1 _09688_ (.A(_04018_),
    .B(_04019_),
    .C(_04028_),
    .D(_04031_),
    .Y(_04033_));
 sg13g2_a21o_1 _09689_ (.A2(_03984_),
    .A1(_03824_),
    .B1(_03800_),
    .X(_04034_));
 sg13g2_nand2_1 _09690_ (.Y(_04035_),
    .A(_03985_),
    .B(_04034_));
 sg13g2_o21ai_1 _09691_ (.B1(_03724_),
    .Y(_04036_),
    .A1(_03726_),
    .A2(_04017_));
 sg13g2_xor2_1 _09692_ (.B(_04036_),
    .A(_03716_),
    .X(_04037_));
 sg13g2_and4_1 _09693_ (.A(_04030_),
    .B(_04033_),
    .C(_04035_),
    .D(_04037_),
    .X(_04038_));
 sg13g2_xnor2_1 _09694_ (.Y(_04039_),
    .A(_03914_),
    .B(_03940_));
 sg13g2_nor2b_1 _09695_ (.A(_03885_),
    .B_N(_03977_),
    .Y(_04040_));
 sg13g2_xnor2_1 _09696_ (.Y(_04041_),
    .A(_03861_),
    .B(_04040_));
 sg13g2_nand4_1 _09697_ (.B(_04038_),
    .C(_04039_),
    .A(_04015_),
    .Y(_04042_),
    .D(_04041_));
 sg13g2_nand3_1 _09698_ (.B(_03828_),
    .C(_03986_),
    .A(_03792_),
    .Y(_04043_));
 sg13g2_nor2b_2 _09699_ (.A(_03987_),
    .B_N(_04043_),
    .Y(_04044_));
 sg13g2_xnor2_1 _09700_ (.Y(_04045_),
    .A(_03935_),
    .B(_03993_));
 sg13g2_xor2_1 _09701_ (.B(_03993_),
    .A(_03935_),
    .X(_04046_));
 sg13g2_o21ai_1 _09702_ (.B1(_03961_),
    .Y(_04047_),
    .A1(_03947_),
    .A2(_03962_));
 sg13g2_xnor2_1 _09703_ (.Y(_04048_),
    .A(_03955_),
    .B(_04047_));
 sg13g2_xor2_1 _09704_ (.B(_04047_),
    .A(_03955_),
    .X(_04049_));
 sg13g2_nor2_1 _09705_ (.A(_03791_),
    .B(_03987_),
    .Y(_04050_));
 sg13g2_xnor2_1 _09706_ (.Y(_04051_),
    .A(_03785_),
    .B(_04050_));
 sg13g2_and3_1 _09707_ (.X(_04052_),
    .A(_03983_),
    .B(_04011_),
    .C(_04013_));
 sg13g2_a21oi_1 _09708_ (.A1(_04006_),
    .A2(_04007_),
    .Y(_04053_),
    .B1(_04044_));
 sg13g2_and4_1 _09709_ (.A(_04005_),
    .B(_04009_),
    .C(_04051_),
    .D(_04053_),
    .X(_04054_));
 sg13g2_nor3_1 _09710_ (.A(_03991_),
    .B(_03995_),
    .C(_04014_),
    .Y(_04055_));
 sg13g2_nor4_1 _09711_ (.A(_04012_),
    .B(_04042_),
    .C(_04046_),
    .D(_04049_),
    .Y(_04056_));
 sg13g2_and4_1 _09712_ (.A(_03990_),
    .B(_04054_),
    .C(_04055_),
    .D(_04056_),
    .X(_04057_));
 sg13g2_nand3_1 _09713_ (.B(_04052_),
    .C(_04057_),
    .A(\cpu.IR[12] ),
    .Y(_04058_));
 sg13g2_a21o_1 _09714_ (.A2(_04057_),
    .A1(_04052_),
    .B1(\cpu.IR[12] ),
    .X(_04059_));
 sg13g2_and3_1 _09715_ (.X(_04060_),
    .A(net3624),
    .B(_04058_),
    .C(_04059_));
 sg13g2_o21ai_1 _09716_ (.B1(_02435_),
    .Y(_04061_),
    .A1(\cpu.IR[14] ),
    .A2(_04060_));
 sg13g2_a21o_1 _09717_ (.A2(_03976_),
    .A1(\cpu.IR[14] ),
    .B1(_04061_),
    .X(_04062_));
 sg13g2_nand2b_1 _09718_ (.Y(_04063_),
    .B(\cpu.IR[3] ),
    .A_N(_00546_));
 sg13g2_nor4_1 _09719_ (.A(\cpu.IR[4] ),
    .B(_02428_),
    .C(_02434_),
    .D(_04063_),
    .Y(_04064_));
 sg13g2_or2_1 _09720_ (.X(_04065_),
    .B(net3415),
    .A(net3423));
 sg13g2_nor2b_1 _09721_ (.A(net3383),
    .B_N(net3116),
    .Y(_04066_));
 sg13g2_nand2b_1 _09722_ (.Y(_04067_),
    .B(net3116),
    .A_N(net3384));
 sg13g2_or4_2 _09723_ (.A(_01696_),
    .B(_01755_),
    .C(_01756_),
    .D(_02434_),
    .X(_04068_));
 sg13g2_nand2_2 _09724_ (.Y(_04069_),
    .A(_00552_),
    .B(_02509_));
 sg13g2_nor2_1 _09725_ (.A(_04068_),
    .B(_04069_),
    .Y(_04070_));
 sg13g2_nor3_2 _09726_ (.A(\cpu.IR[21] ),
    .B(_04068_),
    .C(_04069_),
    .Y(_04071_));
 sg13g2_nor2_1 _09727_ (.A(\cpu.q0 ),
    .B(_04071_),
    .Y(_04072_));
 sg13g2_o21ai_1 _09728_ (.B1(net3406),
    .Y(_04073_),
    .A1(net3635),
    .A2(_04072_));
 sg13g2_nand2_2 _09729_ (.Y(_04074_),
    .A(\cpu.IR[21] ),
    .B(_04070_));
 sg13g2_inv_2 _09730_ (.Y(_04075_),
    .A(_04074_));
 sg13g2_nor3_1 _09731_ (.A(net3107),
    .B(_04073_),
    .C(_04075_),
    .Y(_00013_));
 sg13g2_or3_2 _09732_ (.A(net3918),
    .B(_02424_),
    .C(_02522_),
    .X(cclk));
 sg13g2_a22oi_1 _09733_ (.Y(_04076_),
    .B1(\irqen[4] ),
    .B2(_03505_),
    .A2(\irqen[3] ),
    .A1(net3627));
 sg13g2_nor2b_1 _09734_ (.A(_04071_),
    .B_N(_04076_),
    .Y(_04077_));
 sg13g2_nand2b_1 _09735_ (.Y(_04078_),
    .B(_04076_),
    .A_N(_04071_));
 sg13g2_a22oi_1 _09736_ (.Y(_04079_),
    .B1(_02425_),
    .B2(\irqen[1] ),
    .A2(\irqen[0] ),
    .A1(\uart0.rxvalid ));
 sg13g2_nand2_1 _09737_ (.Y(_04080_),
    .A(\irqen[2] ),
    .B(pwmirq));
 sg13g2_nand3_1 _09738_ (.B(_04079_),
    .C(_04080_),
    .A(net3324),
    .Y(_04081_));
 sg13g2_nor2_1 _09739_ (.A(_04074_),
    .B(_04081_),
    .Y(_04082_));
 sg13g2_a21oi_1 _09740_ (.A1(net3626),
    .A2(_04072_),
    .Y(_00012_),
    .B1(_04082_));
 sg13g2_a21o_1 _09741_ (.A2(_04074_),
    .A1(\cpu.q0 ),
    .B1(_04081_),
    .X(_00014_));
 sg13g2_xor2_1 _09742_ (.B(\tcount[1] ),
    .A(\tcount[0] ),
    .X(_00038_));
 sg13g2_nand3_1 _09743_ (.B(\tcount[1] ),
    .C(\tcount[2] ),
    .A(\tcount[0] ),
    .Y(_04083_));
 sg13g2_a21o_1 _09744_ (.A2(\tcount[1] ),
    .A1(\tcount[0] ),
    .B1(\tcount[2] ),
    .X(_04084_));
 sg13g2_and2_1 _09745_ (.A(_04083_),
    .B(_04084_),
    .X(_00049_));
 sg13g2_nor2_1 _09746_ (.A(_01735_),
    .B(_04083_),
    .Y(_04085_));
 sg13g2_xnor2_1 _09747_ (.Y(_00052_),
    .A(\tcount[3] ),
    .B(_04083_));
 sg13g2_and2_1 _09748_ (.A(\tcount[4] ),
    .B(_04085_),
    .X(_04086_));
 sg13g2_xor2_1 _09749_ (.B(_04085_),
    .A(\tcount[4] ),
    .X(_00053_));
 sg13g2_xor2_1 _09750_ (.B(_04086_),
    .A(\tcount[5] ),
    .X(_00054_));
 sg13g2_nand3_1 _09751_ (.B(\tcount[6] ),
    .C(_04086_),
    .A(\tcount[5] ),
    .Y(_04087_));
 sg13g2_a21o_1 _09752_ (.A2(_04086_),
    .A1(\tcount[5] ),
    .B1(\tcount[6] ),
    .X(_04088_));
 sg13g2_and2_1 _09753_ (.A(_04087_),
    .B(_04088_),
    .X(_00055_));
 sg13g2_nor2_1 _09754_ (.A(_01737_),
    .B(_04087_),
    .Y(_04089_));
 sg13g2_xnor2_1 _09755_ (.Y(_00056_),
    .A(\tcount[7] ),
    .B(_04087_));
 sg13g2_xor2_1 _09756_ (.B(_04089_),
    .A(\tcount[8] ),
    .X(_00057_));
 sg13g2_nand3_1 _09757_ (.B(\tcount[9] ),
    .C(_04089_),
    .A(\tcount[8] ),
    .Y(_04090_));
 sg13g2_a21o_1 _09758_ (.A2(_04089_),
    .A1(\tcount[8] ),
    .B1(\tcount[9] ),
    .X(_04091_));
 sg13g2_and2_1 _09759_ (.A(_04090_),
    .B(_04091_),
    .X(_00058_));
 sg13g2_nor2_1 _09760_ (.A(_01739_),
    .B(_04090_),
    .Y(_04092_));
 sg13g2_xnor2_1 _09761_ (.Y(_00028_),
    .A(\tcount[10] ),
    .B(_04090_));
 sg13g2_xor2_1 _09762_ (.B(_04092_),
    .A(\tcount[11] ),
    .X(_00029_));
 sg13g2_nand3_1 _09763_ (.B(\tcount[12] ),
    .C(_04092_),
    .A(\tcount[11] ),
    .Y(_04093_));
 sg13g2_a21o_1 _09764_ (.A2(_04092_),
    .A1(\tcount[11] ),
    .B1(\tcount[12] ),
    .X(_04094_));
 sg13g2_and2_1 _09765_ (.A(_04093_),
    .B(_04094_),
    .X(_00030_));
 sg13g2_nor2_1 _09766_ (.A(_01740_),
    .B(_04093_),
    .Y(_04095_));
 sg13g2_xnor2_1 _09767_ (.Y(_00031_),
    .A(\tcount[13] ),
    .B(_04093_));
 sg13g2_and2_1 _09768_ (.A(\tcount[14] ),
    .B(_04095_),
    .X(_04096_));
 sg13g2_xor2_1 _09769_ (.B(_04095_),
    .A(\tcount[14] ),
    .X(_00032_));
 sg13g2_xor2_1 _09770_ (.B(_04096_),
    .A(\tcount[15] ),
    .X(_00033_));
 sg13g2_and3_1 _09771_ (.X(_04097_),
    .A(\tcount[16] ),
    .B(\tcount[15] ),
    .C(_04096_));
 sg13g2_a21oi_1 _09772_ (.A1(\tcount[15] ),
    .A2(_04096_),
    .Y(_04098_),
    .B1(\tcount[16] ));
 sg13g2_nor2_1 _09773_ (.A(_04097_),
    .B(_04098_),
    .Y(_00034_));
 sg13g2_xor2_1 _09774_ (.B(_04097_),
    .A(\tcount[17] ),
    .X(_00035_));
 sg13g2_nand3_1 _09775_ (.B(\tcount[18] ),
    .C(_04097_),
    .A(\tcount[17] ),
    .Y(_04099_));
 sg13g2_a21o_1 _09776_ (.A2(_04097_),
    .A1(\tcount[17] ),
    .B1(\tcount[18] ),
    .X(_04100_));
 sg13g2_and2_1 _09777_ (.A(_04099_),
    .B(_04100_),
    .X(_00036_));
 sg13g2_nor2_1 _09778_ (.A(_01736_),
    .B(_04099_),
    .Y(_04101_));
 sg13g2_xnor2_1 _09779_ (.Y(_00037_),
    .A(\tcount[19] ),
    .B(_04099_));
 sg13g2_and2_1 _09780_ (.A(\tcount[20] ),
    .B(_04101_),
    .X(_04102_));
 sg13g2_xor2_1 _09781_ (.B(_04101_),
    .A(\tcount[20] ),
    .X(_00039_));
 sg13g2_xor2_1 _09782_ (.B(_04102_),
    .A(\tcount[21] ),
    .X(_00040_));
 sg13g2_and3_1 _09783_ (.X(_04103_),
    .A(\tcount[21] ),
    .B(\tcount[22] ),
    .C(_04102_));
 sg13g2_a21oi_1 _09784_ (.A1(\tcount[21] ),
    .A2(_04102_),
    .Y(_04104_),
    .B1(\tcount[22] ));
 sg13g2_nor2_1 _09785_ (.A(_04103_),
    .B(_04104_),
    .Y(_00041_));
 sg13g2_xor2_1 _09786_ (.B(_04103_),
    .A(\tcount[23] ),
    .X(_00042_));
 sg13g2_nand3_1 _09787_ (.B(\tcount[24] ),
    .C(_04103_),
    .A(\tcount[23] ),
    .Y(_04105_));
 sg13g2_a21o_1 _09788_ (.A2(_04103_),
    .A1(\tcount[23] ),
    .B1(\tcount[24] ),
    .X(_04106_));
 sg13g2_and2_1 _09789_ (.A(_04105_),
    .B(_04106_),
    .X(_00043_));
 sg13g2_nor2_1 _09790_ (.A(_01738_),
    .B(_04105_),
    .Y(_04107_));
 sg13g2_xnor2_1 _09791_ (.Y(_00044_),
    .A(\tcount[25] ),
    .B(_04105_));
 sg13g2_and2_1 _09792_ (.A(\tcount[26] ),
    .B(_04107_),
    .X(_04108_));
 sg13g2_xor2_1 _09793_ (.B(_04107_),
    .A(\tcount[26] ),
    .X(_00045_));
 sg13g2_xor2_1 _09794_ (.B(_04108_),
    .A(\tcount[27] ),
    .X(_00046_));
 sg13g2_and3_1 _09795_ (.X(_04109_),
    .A(\tcount[27] ),
    .B(\tcount[28] ),
    .C(_04108_));
 sg13g2_a21oi_1 _09796_ (.A1(\tcount[27] ),
    .A2(_04108_),
    .Y(_04110_),
    .B1(\tcount[28] ));
 sg13g2_nor2_1 _09797_ (.A(_04109_),
    .B(_04110_),
    .Y(_00047_));
 sg13g2_xor2_1 _09798_ (.B(_04109_),
    .A(\tcount[29] ),
    .X(_00048_));
 sg13g2_nand3_1 _09799_ (.B(\tcount[30] ),
    .C(_04109_),
    .A(\tcount[29] ),
    .Y(_04111_));
 sg13g2_a21o_1 _09800_ (.A2(_04109_),
    .A1(\tcount[29] ),
    .B1(\tcount[30] ),
    .X(_04112_));
 sg13g2_and2_1 _09801_ (.A(_04111_),
    .B(_04112_),
    .X(_00050_));
 sg13g2_xnor2_1 _09802_ (.Y(_00051_),
    .A(\tcount[31] ),
    .B(_04111_));
 sg13g2_nor3_2 _09803_ (.A(\cpu.Bimm[1] ),
    .B(_01690_),
    .C(_01695_),
    .Y(_04113_));
 sg13g2_nor2_1 _09804_ (.A(net3438),
    .B(_02436_),
    .Y(_04114_));
 sg13g2_nand2_2 _09805_ (.Y(_04115_),
    .A(net3395),
    .B(_02437_));
 sg13g2_nor4_1 _09806_ (.A(\cpu.Bimm[7] ),
    .B(_01651_),
    .C(\cpu.Bimm[5] ),
    .D(\cpu.IR[24] ),
    .Y(_04116_));
 sg13g2_nor2_1 _09807_ (.A(net3644),
    .B(\cpu.Bimm[10] ),
    .Y(_04117_));
 sg13g2_nand4_1 _09808_ (.B(\cpu.Bimm[8] ),
    .C(_04116_),
    .A(\cpu.Bimm[9] ),
    .Y(_04118_),
    .D(_04117_));
 sg13g2_nor4_1 _09809_ (.A(\cpu.IR[23] ),
    .B(\cpu.IR[22] ),
    .C(net3694),
    .D(_02514_),
    .Y(_04119_));
 sg13g2_nand3b_1 _09810_ (.B(net3645),
    .C(_04119_),
    .Y(_04120_),
    .A_N(\cpu.IR[21] ));
 sg13g2_nor3_1 _09811_ (.A(_04068_),
    .B(_04118_),
    .C(_04120_),
    .Y(_04121_));
 sg13g2_nor4_2 _09812_ (.A(net3449),
    .B(net3383),
    .C(net3356),
    .Y(_04122_),
    .D(net3318));
 sg13g2_nand2_2 _09813_ (.Y(_04123_),
    .A(\cpu.Bimm[3] ),
    .B(net3701));
 sg13g2_nor3_2 _09814_ (.A(_01679_),
    .B(_04122_),
    .C(_04123_),
    .Y(_04124_));
 sg13g2_nand2_1 _09815_ (.Y(_04125_),
    .A(_04113_),
    .B(_04124_));
 sg13g2_a21oi_1 _09816_ (.A1(net3699),
    .A2(_03970_),
    .Y(_04126_),
    .B1(_02438_));
 sg13g2_o21ai_1 _09817_ (.B1(_04126_),
    .Y(_04127_),
    .A1(net3699),
    .A2(_03974_));
 sg13g2_nor3_1 _09818_ (.A(net3694),
    .B(_02437_),
    .C(_02514_),
    .Y(_04128_));
 sg13g2_nand3b_1 _09819_ (.B(_02436_),
    .C(_02513_),
    .Y(_04129_),
    .A_N(net3694));
 sg13g2_nor2_1 _09820_ (.A(_03847_),
    .B(net3351),
    .Y(_04130_));
 sg13g2_a21oi_1 _09821_ (.A1(_03778_),
    .A2(net3351),
    .Y(_04131_),
    .B1(_04130_));
 sg13g2_nor2_1 _09822_ (.A(_03729_),
    .B(net3342),
    .Y(_04132_));
 sg13g2_a21oi_1 _09823_ (.A1(_03923_),
    .A2(net3341),
    .Y(_04133_),
    .B1(_04132_));
 sg13g2_nand2_1 _09824_ (.Y(_04134_),
    .A(_03863_),
    .B(net3350));
 sg13g2_a21oi_1 _09825_ (.A1(_03794_),
    .A2(net3342),
    .Y(_04135_),
    .B1(net3265));
 sg13g2_a22oi_1 _09826_ (.Y(_04136_),
    .B1(_04134_),
    .B2(_04135_),
    .A2(_04133_),
    .A1(net3261));
 sg13g2_a21oi_1 _09827_ (.A1(_03686_),
    .A2(net3345),
    .Y(_04137_),
    .B1(net3266));
 sg13g2_o21ai_1 _09828_ (.B1(_04137_),
    .Y(_04138_),
    .A1(_03950_),
    .A2(net3344));
 sg13g2_a21oi_1 _09829_ (.A1(net3262),
    .A2(_04131_),
    .Y(_04139_),
    .B1(net3279));
 sg13g2_a22oi_1 _09830_ (.Y(_04140_),
    .B1(_04138_),
    .B2(_04139_),
    .A2(_04136_),
    .A1(net3280));
 sg13g2_nand2_1 _09831_ (.Y(_04141_),
    .A(net3277),
    .B(_04140_));
 sg13g2_and2_1 _09832_ (.A(_03888_),
    .B(net3342),
    .X(_04142_));
 sg13g2_a21oi_1 _09833_ (.A1(_03819_),
    .A2(net3349),
    .Y(_04143_),
    .B1(_04142_));
 sg13g2_o21ai_1 _09834_ (.B1(net3268),
    .Y(_04144_),
    .A1(_03718_),
    .A2(net3352));
 sg13g2_a21oi_1 _09835_ (.A1(_03930_),
    .A2(net3352),
    .Y(_04145_),
    .B1(_04144_));
 sg13g2_a21oi_1 _09836_ (.A1(net3262),
    .A2(_04143_),
    .Y(_04146_),
    .B1(_04145_));
 sg13g2_nor2_1 _09837_ (.A(net3279),
    .B(_04146_),
    .Y(_04147_));
 sg13g2_nor2_1 _09838_ (.A(_03665_),
    .B(net3351),
    .Y(_04148_));
 sg13g2_a21oi_1 _09839_ (.A1(_02432_),
    .A2(net3349),
    .Y(_04149_),
    .B1(_04148_));
 sg13g2_o21ai_1 _09840_ (.B1(net3268),
    .Y(_04150_),
    .A1(_03854_),
    .A2(net3339));
 sg13g2_a21oi_1 _09841_ (.A1(_03762_),
    .A2(net3341),
    .Y(_04151_),
    .B1(_04150_));
 sg13g2_a21oi_1 _09842_ (.A1(net3264),
    .A2(_04149_),
    .Y(_04152_),
    .B1(_04151_));
 sg13g2_a21oi_1 _09843_ (.A1(net3281),
    .A2(_04152_),
    .Y(_04153_),
    .B1(_04147_));
 sg13g2_o21ai_1 _09844_ (.B1(_04141_),
    .Y(_04154_),
    .A1(net3277),
    .A2(_04153_));
 sg13g2_nand2_1 _09845_ (.Y(_04155_),
    .A(_03880_),
    .B(net3339));
 sg13g2_o21ai_1 _09846_ (.B1(_04155_),
    .Y(_04156_),
    .A1(_03769_),
    .A2(net3339));
 sg13g2_nand2_1 _09847_ (.Y(_04157_),
    .A(_03936_),
    .B(net3346));
 sg13g2_o21ai_1 _09848_ (.B1(_04157_),
    .Y(_04158_),
    .A1(_03707_),
    .A2(net3345));
 sg13g2_nand2_1 _09849_ (.Y(_04159_),
    .A(_03896_),
    .B(net3352));
 sg13g2_a21oi_1 _09850_ (.A1(_03812_),
    .A2(net3345),
    .Y(_04160_),
    .B1(net3267));
 sg13g2_a22oi_1 _09851_ (.Y(_04161_),
    .B1(_04159_),
    .B2(_04160_),
    .A2(_04158_),
    .A1(net3267));
 sg13g2_a21o_1 _09852_ (.A2(net3354),
    .A1(_03657_),
    .B1(net3266),
    .X(_04162_));
 sg13g2_a21oi_1 _09853_ (.A1(_02501_),
    .A2(net3345),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_o21ai_1 _09854_ (.B1(net3288),
    .Y(_04164_),
    .A1(net3269),
    .A2(_04156_));
 sg13g2_o21ai_1 _09855_ (.B1(net3277),
    .Y(_04165_),
    .A1(_04163_),
    .A2(_04164_));
 sg13g2_a21oi_1 _09856_ (.A1(net3284),
    .A2(_04161_),
    .Y(_04166_),
    .B1(_04165_));
 sg13g2_a21oi_1 _09857_ (.A1(_03739_),
    .A2(net3344),
    .Y(_04167_),
    .B1(net3265));
 sg13g2_o21ai_1 _09858_ (.B1(_04167_),
    .Y(_04168_),
    .A1(_03916_),
    .A2(net3344));
 sg13g2_nand2_1 _09859_ (.Y(_04169_),
    .A(_03871_),
    .B(net3342));
 sg13g2_o21ai_1 _09860_ (.B1(_04169_),
    .Y(_04170_),
    .A1(_03803_),
    .A2(net3344));
 sg13g2_o21ai_1 _09861_ (.B1(_04168_),
    .Y(_04171_),
    .A1(net3269),
    .A2(_04170_));
 sg13g2_nor2_1 _09862_ (.A(_03957_),
    .B(net3349),
    .Y(_04172_));
 sg13g2_a21oi_1 _09863_ (.A1(_03675_),
    .A2(net3349),
    .Y(_04173_),
    .B1(_04172_));
 sg13g2_nand2_1 _09864_ (.Y(_04174_),
    .A(_03837_),
    .B(net3351));
 sg13g2_a21oi_1 _09865_ (.A1(_03786_),
    .A2(net3341),
    .Y(_04175_),
    .B1(net3261));
 sg13g2_a22oi_1 _09866_ (.Y(_04176_),
    .B1(_04174_),
    .B2(_04175_),
    .A2(_04173_),
    .A1(net3261));
 sg13g2_nand2_1 _09867_ (.Y(_04177_),
    .A(net3280),
    .B(_04176_));
 sg13g2_o21ai_1 _09868_ (.B1(_04177_),
    .Y(_04178_),
    .A1(net3280),
    .A2(_04171_));
 sg13g2_a21oi_1 _09869_ (.A1(net3273),
    .A2(_04178_),
    .Y(_04179_),
    .B1(_04166_));
 sg13g2_mux2_1 _09870_ (.A0(_04154_),
    .A1(_04179_),
    .S(net3304),
    .X(_04180_));
 sg13g2_nand2_1 _09871_ (.Y(_04181_),
    .A(_03854_),
    .B(net3339));
 sg13g2_o21ai_1 _09872_ (.B1(_04181_),
    .Y(_04182_),
    .A1(_03762_),
    .A2(net3341));
 sg13g2_o21ai_1 _09873_ (.B1(net3268),
    .Y(_04183_),
    .A1(_02432_),
    .A2(net3349));
 sg13g2_a21oi_1 _09874_ (.A1(_03665_),
    .A2(net3350),
    .Y(_04184_),
    .B1(_04183_));
 sg13g2_o21ai_1 _09875_ (.B1(net3287),
    .Y(_04185_),
    .A1(net3269),
    .A2(_04182_));
 sg13g2_nor2_1 _09876_ (.A(_03718_),
    .B(net3344),
    .Y(_04186_));
 sg13g2_a21oi_1 _09877_ (.A1(_03930_),
    .A2(net3346),
    .Y(_04187_),
    .B1(_04186_));
 sg13g2_nand2_1 _09878_ (.Y(_04188_),
    .A(_03888_),
    .B(net3350));
 sg13g2_a21oi_1 _09879_ (.A1(_03819_),
    .A2(net3341),
    .Y(_04189_),
    .B1(net3262));
 sg13g2_a22oi_1 _09880_ (.Y(_04190_),
    .B1(_04188_),
    .B2(_04189_),
    .A2(_04187_),
    .A1(net3261));
 sg13g2_a21oi_1 _09881_ (.A1(_03923_),
    .A2(net3349),
    .Y(_04191_),
    .B1(net3265));
 sg13g2_o21ai_1 _09882_ (.B1(_04191_),
    .Y(_04192_),
    .A1(_03729_),
    .A2(net3349));
 sg13g2_and2_1 _09883_ (.A(_03794_),
    .B(net3350),
    .X(_04193_));
 sg13g2_a21oi_1 _09884_ (.A1(_03863_),
    .A2(net3341),
    .Y(_04194_),
    .B1(_04193_));
 sg13g2_a21oi_1 _09885_ (.A1(net3261),
    .A2(_04194_),
    .Y(_04195_),
    .B1(net3279));
 sg13g2_nor2_1 _09886_ (.A(_03949_),
    .B(net3348),
    .Y(_04196_));
 sg13g2_a21oi_2 _09887_ (.B1(_04196_),
    .Y(_04197_),
    .A2(net3348),
    .A1(_03687_));
 sg13g2_a21oi_1 _09888_ (.A1(_03778_),
    .A2(net3339),
    .Y(_04198_),
    .B1(net3261));
 sg13g2_o21ai_1 _09889_ (.B1(_04198_),
    .Y(_04199_),
    .A1(_03847_),
    .A2(net3340));
 sg13g2_o21ai_1 _09890_ (.B1(_04199_),
    .Y(_04200_),
    .A1(net3268),
    .A2(_04197_));
 sg13g2_nor2_1 _09891_ (.A(net3287),
    .B(_04200_),
    .Y(_04201_));
 sg13g2_a21oi_1 _09892_ (.A1(_04192_),
    .A2(_04195_),
    .Y(_04202_),
    .B1(_04201_));
 sg13g2_o21ai_1 _09893_ (.B1(net3276),
    .Y(_04203_),
    .A1(_04184_),
    .A2(_04185_));
 sg13g2_a21oi_1 _09894_ (.A1(net3279),
    .A2(_04190_),
    .Y(_04204_),
    .B1(_04203_));
 sg13g2_a21oi_1 _09895_ (.A1(net3270),
    .A2(_04202_),
    .Y(_04205_),
    .B1(_04204_));
 sg13g2_nand2_1 _09896_ (.Y(_04206_),
    .A(_03916_),
    .B(net3344));
 sg13g2_o21ai_1 _09897_ (.B1(_04206_),
    .Y(_04207_),
    .A1(_03739_),
    .A2(net3344));
 sg13g2_nand2_1 _09898_ (.Y(_04208_),
    .A(_03802_),
    .B(net3342));
 sg13g2_a21oi_1 _09899_ (.A1(_03871_),
    .A2(net3349),
    .Y(_04209_),
    .B1(net3265));
 sg13g2_a22oi_1 _09900_ (.Y(_04210_),
    .B1(_04208_),
    .B2(_04209_),
    .A2(_04207_),
    .A1(net3265));
 sg13g2_o21ai_1 _09901_ (.B1(net3268),
    .Y(_04211_),
    .A1(_03957_),
    .A2(net3342));
 sg13g2_a21o_1 _09902_ (.A2(net3341),
    .A1(_03675_),
    .B1(_04211_),
    .X(_04212_));
 sg13g2_and2_1 _09903_ (.A(_03837_),
    .B(net3339),
    .X(_04213_));
 sg13g2_a21oi_1 _09904_ (.A1(_03786_),
    .A2(net3351),
    .Y(_04214_),
    .B1(_04213_));
 sg13g2_a21oi_1 _09905_ (.A1(net3262),
    .A2(_04214_),
    .Y(_04215_),
    .B1(net3279));
 sg13g2_mux2_1 _09906_ (.A0(_03812_),
    .A1(_03896_),
    .S(net3346),
    .X(_04216_));
 sg13g2_nand2_1 _09907_ (.Y(_04217_),
    .A(_03936_),
    .B(net3352));
 sg13g2_a21oi_1 _09908_ (.A1(_03706_),
    .A2(net3345),
    .Y(_04218_),
    .B1(net3266));
 sg13g2_a221oi_1 _09909_ (.B2(_04218_),
    .C1(net3279),
    .B1(_04217_),
    .A1(net3266),
    .Y(_04219_),
    .A2(_04216_));
 sg13g2_nand2_1 _09910_ (.Y(_04220_),
    .A(_03879_),
    .B(net3351));
 sg13g2_a21oi_1 _09911_ (.A1(_03769_),
    .A2(net3341),
    .Y(_04221_),
    .B1(net3262));
 sg13g2_nand2_1 _09912_ (.Y(_04222_),
    .A(_03657_),
    .B(net3345));
 sg13g2_o21ai_1 _09913_ (.B1(_04222_),
    .Y(_04223_),
    .A1(_02502_),
    .A2(net3345));
 sg13g2_a22oi_1 _09914_ (.Y(_04224_),
    .B1(_04223_),
    .B2(net3262),
    .A2(_04221_),
    .A1(_04220_));
 sg13g2_a21oi_1 _09915_ (.A1(net3280),
    .A2(_04224_),
    .Y(_04225_),
    .B1(_04219_));
 sg13g2_a221oi_1 _09916_ (.B2(_04215_),
    .C1(net3270),
    .B1(_04212_),
    .A1(net3279),
    .Y(_04226_),
    .A2(_04210_));
 sg13g2_a21o_1 _09917_ (.A2(_04225_),
    .A1(net3270),
    .B1(_04226_),
    .X(_04227_));
 sg13g2_nand2_1 _09918_ (.Y(_04228_),
    .A(net3303),
    .B(_04205_));
 sg13g2_o21ai_1 _09919_ (.B1(_04228_),
    .Y(_04229_),
    .A1(net3304),
    .A2(_04227_));
 sg13g2_nor2_1 _09920_ (.A(net3296),
    .B(_04229_),
    .Y(_04230_));
 sg13g2_a21oi_1 _09921_ (.A1(net3296),
    .A2(_04180_),
    .Y(_04231_),
    .B1(_04230_));
 sg13g2_nand2_1 _09922_ (.Y(_04232_),
    .A(net3347),
    .B(_04231_));
 sg13g2_nor4_2 _09923_ (.A(_00562_),
    .B(_00552_),
    .C(_02437_),
    .Y(_04233_),
    .D(_02514_));
 sg13g2_nor2_1 _09924_ (.A(net3306),
    .B(_04233_),
    .Y(_04234_));
 sg13g2_and2_1 _09925_ (.A(_04223_),
    .B(_04233_),
    .X(_04235_));
 sg13g2_nand2_2 _09926_ (.Y(_04236_),
    .A(_04223_),
    .B(_04233_));
 sg13g2_nand2_2 _09927_ (.Y(_04237_),
    .A(net3272),
    .B(_04236_));
 sg13g2_nor2_2 _09928_ (.A(net3288),
    .B(_04235_),
    .Y(_04238_));
 sg13g2_nand2_1 _09929_ (.Y(_04239_),
    .A(net3284),
    .B(_04236_));
 sg13g2_nor2_2 _09930_ (.A(net3269),
    .B(_04235_),
    .Y(_04240_));
 sg13g2_nand2_1 _09931_ (.Y(_04241_),
    .A(net3266),
    .B(_04236_));
 sg13g2_and2_1 _09932_ (.A(_04223_),
    .B(net3129),
    .X(_04242_));
 sg13g2_nand2_1 _09933_ (.Y(_04243_),
    .A(_04239_),
    .B(_04242_));
 sg13g2_nand2_1 _09934_ (.Y(_04244_),
    .A(net3278),
    .B(_04243_));
 sg13g2_nand2_1 _09935_ (.Y(_04245_),
    .A(_04237_),
    .B(_04244_));
 sg13g2_nor2_1 _09936_ (.A(_04234_),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_o21ai_1 _09937_ (.B1(_04246_),
    .Y(_04247_),
    .A1(net3296),
    .A2(_04233_));
 sg13g2_a21oi_1 _09938_ (.A1(net3353),
    .A2(_04247_),
    .Y(_04248_),
    .B1(_02514_));
 sg13g2_nand2_1 _09939_ (.Y(_04249_),
    .A(net3694),
    .B(net3695));
 sg13g2_nor2_1 _09940_ (.A(net3699),
    .B(_04249_),
    .Y(_04250_));
 sg13g2_nand2b_1 _09941_ (.Y(_04251_),
    .B(_01697_),
    .A_N(_04249_));
 sg13g2_a21o_1 _09942_ (.A2(_02502_),
    .A1(net3289),
    .B1(net3409),
    .X(_04252_));
 sg13g2_nor2_2 _09943_ (.A(_01697_),
    .B(_04249_),
    .Y(_04253_));
 sg13g2_nand3_1 _09944_ (.B(net3699),
    .C(net3695),
    .A(net3694),
    .Y(_04254_));
 sg13g2_nand3b_1 _09945_ (.B(_02501_),
    .C(_04253_),
    .Y(_04255_),
    .A_N(net3289));
 sg13g2_nand4_1 _09946_ (.B(_04127_),
    .C(_04252_),
    .A(_02512_),
    .Y(_04256_),
    .D(_04255_));
 sg13g2_a21oi_1 _09947_ (.A1(_04232_),
    .A2(_04248_),
    .Y(_04257_),
    .B1(_04256_));
 sg13g2_a21oi_1 _09948_ (.A1(_02505_),
    .A2(_03567_),
    .Y(_04258_),
    .B1(_02512_));
 sg13g2_o21ai_1 _09949_ (.B1(_04258_),
    .Y(_04259_),
    .A1(_02505_),
    .A2(\cdi[24] ));
 sg13g2_a21oi_2 _09950_ (.B1(_02507_),
    .Y(_04260_),
    .A2(net3236),
    .A1(_01697_));
 sg13g2_a22oi_1 _09951_ (.Y(_04261_),
    .B1(\cdi[16] ),
    .B2(_04260_),
    .A2(\cdi[0] ),
    .A1(_02517_));
 sg13g2_a21o_1 _09952_ (.A2(_04261_),
    .A1(_04259_),
    .B1(_01764_),
    .X(_04262_));
 sg13g2_o21ai_1 _09953_ (.B1(_04262_),
    .Y(_04263_),
    .A1(net3358),
    .A2(_04257_));
 sg13g2_mux2_1 _09954_ (.A0(net3047),
    .A1(\cpu.regs[13][0] ),
    .S(net3220),
    .X(_00695_));
 sg13g2_nor2_1 _09955_ (.A(_02514_),
    .B(net3353),
    .Y(_04264_));
 sg13g2_nand2_1 _09956_ (.Y(_04265_),
    .A(_02513_),
    .B(net3347));
 sg13g2_nand2_1 _09957_ (.Y(_04266_),
    .A(net3304),
    .B(_04154_));
 sg13g2_nand2_1 _09958_ (.Y(_04267_),
    .A(net3288),
    .B(_04161_));
 sg13g2_o21ai_1 _09959_ (.B1(_04241_),
    .Y(_04268_),
    .A1(net3266),
    .A2(_04156_));
 sg13g2_o21ai_1 _09960_ (.B1(_04267_),
    .Y(_04269_),
    .A1(net3288),
    .A2(_04268_));
 sg13g2_nand2_1 _09961_ (.Y(_04270_),
    .A(net3277),
    .B(_04178_));
 sg13g2_o21ai_1 _09962_ (.B1(_04270_),
    .Y(_04271_),
    .A1(net3277),
    .A2(_04269_));
 sg13g2_o21ai_1 _09963_ (.B1(_04266_),
    .Y(_04272_),
    .A1(net3304),
    .A2(_04271_));
 sg13g2_nand2_1 _09964_ (.Y(_04273_),
    .A(net3296),
    .B(_04229_));
 sg13g2_o21ai_1 _09965_ (.B1(_04273_),
    .Y(_04274_),
    .A1(net3296),
    .A2(_04272_));
 sg13g2_nor2_1 _09966_ (.A(net3311),
    .B(_04274_),
    .Y(_04275_));
 sg13g2_a21o_1 _09967_ (.A2(_04149_),
    .A1(net3268),
    .B1(_04240_),
    .X(_04276_));
 sg13g2_a21oi_1 _09968_ (.A1(net3285),
    .A2(_04276_),
    .Y(_04277_),
    .B1(_04238_));
 sg13g2_o21ai_1 _09969_ (.B1(_04237_),
    .Y(_04278_),
    .A1(net3272),
    .A2(_04277_));
 sg13g2_a21oi_1 _09970_ (.A1(_04237_),
    .A2(_04244_),
    .Y(_04279_),
    .B1(net3306));
 sg13g2_a21oi_1 _09971_ (.A1(net3306),
    .A2(_04278_),
    .Y(_04280_),
    .B1(_04234_));
 sg13g2_nor2b_1 _09972_ (.A(_04279_),
    .B_N(_04280_),
    .Y(_04281_));
 sg13g2_mux2_2 _09973_ (.A0(_04246_),
    .A1(_04281_),
    .S(net3295),
    .X(_04282_));
 sg13g2_nand2_1 _09974_ (.Y(_04283_),
    .A(net3353),
    .B(_04282_));
 sg13g2_nor2b_1 _09975_ (.A(net3438),
    .B_N(_04069_),
    .Y(_04284_));
 sg13g2_nand2_1 _09976_ (.Y(_04285_),
    .A(net3393),
    .B(_04069_));
 sg13g2_nor2_1 _09977_ (.A(_02433_),
    .B(net3304),
    .Y(_04286_));
 sg13g2_nor2_1 _09978_ (.A(_00552_),
    .B(_02510_),
    .Y(_04287_));
 sg13g2_o21ai_1 _09979_ (.B1(net3375),
    .Y(_04288_),
    .A1(_02433_),
    .A2(net3304));
 sg13g2_a22oi_1 _09980_ (.Y(_04289_),
    .B1(net3409),
    .B2(_04288_),
    .A2(net3304),
    .A1(_02433_));
 sg13g2_a221oi_1 _09981_ (.B2(_04253_),
    .C1(_04289_),
    .B1(_04286_),
    .A1(net3140),
    .Y(_04290_),
    .A2(net3338));
 sg13g2_nand2_1 _09982_ (.Y(_04291_),
    .A(_04283_),
    .B(_04290_));
 sg13g2_o21ai_1 _09983_ (.B1(_04115_),
    .Y(_04292_),
    .A1(_04275_),
    .A2(_04291_));
 sg13g2_nand2_1 _09984_ (.Y(_04293_),
    .A(net3134),
    .B(\cdi[9] ));
 sg13g2_o21ai_1 _09985_ (.B1(_04293_),
    .Y(_04294_),
    .A1(net3134),
    .A2(_03581_));
 sg13g2_o21ai_1 _09986_ (.B1(net3448),
    .Y(_04295_),
    .A1(_02518_),
    .A2(\cdi[1] ));
 sg13g2_a21oi_1 _09987_ (.A1(_03476_),
    .A2(_04260_),
    .Y(_04296_),
    .B1(_04295_));
 sg13g2_o21ai_1 _09988_ (.B1(_04296_),
    .Y(_04297_),
    .A1(_02512_),
    .A2(_04294_));
 sg13g2_nand2_1 _09989_ (.Y(_04298_),
    .A(_04292_),
    .B(_04297_));
 sg13g2_mux2_1 _09990_ (.A0(net3042),
    .A1(\cpu.regs[13][1] ),
    .S(net3225),
    .X(_00696_));
 sg13g2_mux2_1 _09991_ (.A0(\cdi[10] ),
    .A1(\cdi[26] ),
    .S(net3140),
    .X(_04299_));
 sg13g2_o21ai_1 _09992_ (.B1(net3448),
    .Y(_04300_),
    .A1(_02518_),
    .A2(\cdi[2] ));
 sg13g2_a21oi_1 _09993_ (.A1(_03493_),
    .A2(_04260_),
    .Y(_04301_),
    .B1(_04300_));
 sg13g2_o21ai_1 _09994_ (.B1(_04301_),
    .Y(_04302_),
    .A1(_02512_),
    .A2(_04299_));
 sg13g2_a21oi_1 _09995_ (.A1(net3268),
    .A2(_04197_),
    .Y(_04303_),
    .B1(_04240_));
 sg13g2_inv_1 _09996_ (.Y(_04304_),
    .A(_04303_));
 sg13g2_a21oi_2 _09997_ (.B1(_04238_),
    .Y(_04305_),
    .A2(_04304_),
    .A1(net3286));
 sg13g2_o21ai_1 _09998_ (.B1(_04237_),
    .Y(_04306_),
    .A1(net3272),
    .A2(_04305_));
 sg13g2_a21oi_1 _09999_ (.A1(net3306),
    .A2(_04306_),
    .Y(_04307_),
    .B1(_04279_));
 sg13g2_mux2_1 _10000_ (.A0(_04281_),
    .A1(_04307_),
    .S(net3297),
    .X(_04308_));
 sg13g2_a21oi_1 _10001_ (.A1(net3269),
    .A2(_04182_),
    .Y(_04309_),
    .B1(_04240_));
 sg13g2_nand2_1 _10002_ (.Y(_04310_),
    .A(net3287),
    .B(_04190_));
 sg13g2_o21ai_1 _10003_ (.B1(_04310_),
    .Y(_04311_),
    .A1(net3287),
    .A2(_04309_));
 sg13g2_nor2_1 _10004_ (.A(net3276),
    .B(_04311_),
    .Y(_04312_));
 sg13g2_a21oi_2 _10005_ (.B1(_04312_),
    .Y(_04313_),
    .A2(_04202_),
    .A1(net3276));
 sg13g2_nor2_1 _10006_ (.A(net3303),
    .B(_04313_),
    .Y(_04314_));
 sg13g2_a21oi_1 _10007_ (.A1(net3303),
    .A2(_04227_),
    .Y(_04315_),
    .B1(_04314_));
 sg13g2_nand2_1 _10008_ (.Y(_04316_),
    .A(net3296),
    .B(_04272_));
 sg13g2_o21ai_1 _10009_ (.B1(_04316_),
    .Y(_04317_),
    .A1(net3296),
    .A2(_04315_));
 sg13g2_nand2_1 _10010_ (.Y(_04318_),
    .A(net3313),
    .B(_04317_));
 sg13g2_nand2_1 _10011_ (.Y(_04319_),
    .A(_03687_),
    .B(net3273));
 sg13g2_a21o_1 _10012_ (.A2(_04319_),
    .A1(net3374),
    .B1(net3411),
    .X(_04320_));
 sg13g2_o21ai_1 _10013_ (.B1(_04320_),
    .Y(_04321_),
    .A1(_03687_),
    .A2(net3273));
 sg13g2_o21ai_1 _10014_ (.B1(_04321_),
    .Y(_04322_),
    .A1(net3454),
    .A2(_04319_));
 sg13g2_a221oi_1 _10015_ (.B2(net3353),
    .C1(_04322_),
    .B1(_04308_),
    .A1(_04025_),
    .Y(_04323_),
    .A2(net3338));
 sg13g2_a21oi_2 _10016_ (.B1(net3358),
    .Y(_04324_),
    .A2(_04323_),
    .A1(_04318_));
 sg13g2_a221oi_1 _10017_ (.B2(\cpu.PCreg0[2] ),
    .C1(_04324_),
    .B1(net3317),
    .A1(\cpu.PC[2] ),
    .Y(_04325_),
    .A2(net3383));
 sg13g2_nand2_1 _10018_ (.Y(_04326_),
    .A(_04302_),
    .B(_04325_));
 sg13g2_mux2_1 _10019_ (.A0(net3039),
    .A1(\cpu.regs[13][2] ),
    .S(net3220),
    .X(_00697_));
 sg13g2_mux2_1 _10020_ (.A0(\cdi[11] ),
    .A1(\cdi[27] ),
    .S(net3137),
    .X(_04327_));
 sg13g2_inv_1 _10021_ (.Y(_04328_),
    .A(_04327_));
 sg13g2_o21ai_1 _10022_ (.B1(net3129),
    .Y(_04329_),
    .A1(net3263),
    .A2(_04131_));
 sg13g2_and2_1 _10023_ (.A(net3287),
    .B(_04136_),
    .X(_04330_));
 sg13g2_a21oi_1 _10024_ (.A1(net3281),
    .A2(_04329_),
    .Y(_04331_),
    .B1(_04330_));
 sg13g2_nor2_1 _10025_ (.A(net3276),
    .B(_04331_),
    .Y(_04332_));
 sg13g2_a21oi_1 _10026_ (.A1(net3277),
    .A2(_04153_),
    .Y(_04333_),
    .B1(_04332_));
 sg13g2_nor2_1 _10027_ (.A(net3303),
    .B(_04333_),
    .Y(_04334_));
 sg13g2_a21oi_1 _10028_ (.A1(net3303),
    .A2(_04271_),
    .Y(_04335_),
    .B1(_04334_));
 sg13g2_nand2_1 _10029_ (.Y(_04336_),
    .A(net3296),
    .B(_04315_));
 sg13g2_o21ai_1 _10030_ (.B1(_04336_),
    .Y(_04337_),
    .A1(net3289),
    .A2(_04335_));
 sg13g2_nor2_1 _10031_ (.A(net3311),
    .B(_04337_),
    .Y(_04338_));
 sg13g2_o21ai_1 _10032_ (.B1(net3129),
    .Y(_04339_),
    .A1(net3263),
    .A2(_04173_));
 sg13g2_a21oi_1 _10033_ (.A1(net3285),
    .A2(_04339_),
    .Y(_04340_),
    .B1(_04238_));
 sg13g2_o21ai_1 _10034_ (.B1(_04237_),
    .Y(_04341_),
    .A1(net3272),
    .A2(_04340_));
 sg13g2_mux2_1 _10035_ (.A0(_04278_),
    .A1(_04341_),
    .S(net3306),
    .X(_04342_));
 sg13g2_nand2_1 _10036_ (.Y(_04343_),
    .A(net3295),
    .B(_04342_));
 sg13g2_o21ai_1 _10037_ (.B1(_04343_),
    .Y(_04344_),
    .A1(net3295),
    .A2(_04307_));
 sg13g2_inv_1 _10038_ (.Y(_04345_),
    .A(_04344_));
 sg13g2_nand2_1 _10039_ (.Y(_04346_),
    .A(_03676_),
    .B(net3284));
 sg13g2_nand2_1 _10040_ (.Y(_04347_),
    .A(net3375),
    .B(_04346_));
 sg13g2_a22oi_1 _10041_ (.Y(_04348_),
    .B1(net3409),
    .B2(_04347_),
    .A2(net3288),
    .A1(_03675_));
 sg13g2_a221oi_1 _10042_ (.B2(net3352),
    .C1(_04348_),
    .B1(_04345_),
    .A1(_04023_),
    .Y(_04349_),
    .A2(net3338));
 sg13g2_o21ai_1 _10043_ (.B1(_04349_),
    .Y(_04350_),
    .A1(net3455),
    .A2(_04346_));
 sg13g2_o21ai_1 _10044_ (.B1(_04115_),
    .Y(_04351_),
    .A1(_04338_),
    .A2(_04350_));
 sg13g2_o21ai_1 _10045_ (.B1(net3448),
    .Y(_04352_),
    .A1(_02518_),
    .A2(\cdi[3] ));
 sg13g2_a221oi_1 _10046_ (.B2(_02511_),
    .C1(_04352_),
    .B1(_04328_),
    .A1(_03502_),
    .Y(_04353_),
    .A2(_04260_));
 sg13g2_a221oi_1 _10047_ (.B2(\cpu.PCreg0[3] ),
    .C1(_04353_),
    .B1(net3317),
    .A1(\cpu.PC[3] ),
    .Y(_04354_),
    .A2(net3384));
 sg13g2_nand2_2 _10048_ (.Y(_04355_),
    .A(_04351_),
    .B(_04354_));
 sg13g2_mux2_1 _10049_ (.A0(net3006),
    .A1(\cpu.regs[13][3] ),
    .S(net3222),
    .X(_00698_));
 sg13g2_o21ai_1 _10050_ (.B1(net3235),
    .Y(_04356_),
    .A1(net3138),
    .A2(\cdi[12] ));
 sg13g2_a21oi_1 _10051_ (.A1(net3137),
    .A2(_03595_),
    .Y(_04357_),
    .B1(_04356_));
 sg13g2_nor2_1 _10052_ (.A(net3134),
    .B(_03516_),
    .Y(_04358_));
 sg13g2_a21oi_1 _10053_ (.A1(net3134),
    .A2(\cdi[4] ),
    .Y(_04359_),
    .B1(_04358_));
 sg13g2_o21ai_1 _10054_ (.B1(net3459),
    .Y(_04360_),
    .A1(net3236),
    .A2(_04359_));
 sg13g2_o21ai_1 _10055_ (.B1(net3448),
    .Y(_04361_),
    .A1(net3625),
    .A2(\cdi[4] ));
 sg13g2_a21oi_1 _10056_ (.A1(_02513_),
    .A2(_04359_),
    .Y(_04362_),
    .B1(_04361_));
 sg13g2_o21ai_1 _10057_ (.B1(_04362_),
    .Y(_04363_),
    .A1(_04357_),
    .A2(_04360_));
 sg13g2_o21ai_1 _10058_ (.B1(net3129),
    .Y(_04364_),
    .A1(net3263),
    .A2(_04214_));
 sg13g2_mux2_1 _10059_ (.A0(_04210_),
    .A1(_04364_),
    .S(net3279),
    .X(_04365_));
 sg13g2_nor2_1 _10060_ (.A(net3276),
    .B(_04365_),
    .Y(_04366_));
 sg13g2_a21oi_1 _10061_ (.A1(net3277),
    .A2(_04225_),
    .Y(_04367_),
    .B1(_04366_));
 sg13g2_mux2_1 _10062_ (.A0(_04367_),
    .A1(_04313_),
    .S(net3303),
    .X(_04368_));
 sg13g2_nor2_1 _10063_ (.A(net3289),
    .B(_04368_),
    .Y(_04369_));
 sg13g2_a21oi_2 _10064_ (.B1(_04369_),
    .Y(_04370_),
    .A2(_04335_),
    .A1(net3289));
 sg13g2_nor2_1 _10065_ (.A(net3311),
    .B(_04370_),
    .Y(_04371_));
 sg13g2_o21ai_1 _10066_ (.B1(net3129),
    .Y(_04372_),
    .A1(net3263),
    .A2(_04207_));
 sg13g2_a21oi_1 _10067_ (.A1(net3286),
    .A2(_04372_),
    .Y(_04373_),
    .B1(_04238_));
 sg13g2_nand2_1 _10068_ (.Y(_04374_),
    .A(net3278),
    .B(_04373_));
 sg13g2_o21ai_1 _10069_ (.B1(_04374_),
    .Y(_04375_),
    .A1(net3278),
    .A2(_04243_));
 sg13g2_nand2_1 _10070_ (.Y(_04376_),
    .A(net3305),
    .B(_04375_));
 sg13g2_o21ai_1 _10071_ (.B1(_04376_),
    .Y(_04377_),
    .A1(net3305),
    .A2(_04306_));
 sg13g2_nor2_1 _10072_ (.A(net3295),
    .B(_04342_),
    .Y(_04378_));
 sg13g2_a21oi_2 _10073_ (.B1(_04378_),
    .Y(_04379_),
    .A2(_04377_),
    .A1(net3295));
 sg13g2_nor2_1 _10074_ (.A(_04027_),
    .B(net3378),
    .Y(_04380_));
 sg13g2_nand2_1 _10075_ (.Y(_04381_),
    .A(_03740_),
    .B(net3266));
 sg13g2_nor2_1 _10076_ (.A(net3454),
    .B(_04381_),
    .Y(_04382_));
 sg13g2_nand2_1 _10077_ (.Y(_04383_),
    .A(net3374),
    .B(_04381_));
 sg13g2_a22oi_1 _10078_ (.Y(_04384_),
    .B1(net3409),
    .B2(_04383_),
    .A2(net3269),
    .A1(_03739_));
 sg13g2_nor3_1 _10079_ (.A(_04380_),
    .B(_04382_),
    .C(_04384_),
    .Y(_04385_));
 sg13g2_o21ai_1 _10080_ (.B1(_04385_),
    .Y(_04386_),
    .A1(net3347),
    .A2(_04379_));
 sg13g2_o21ai_1 _10081_ (.B1(net3356),
    .Y(_04387_),
    .A1(_04371_),
    .A2(_04386_));
 sg13g2_a22oi_1 _10082_ (.Y(_04388_),
    .B1(net3317),
    .B2(\cpu.PCreg0[4] ),
    .A2(net3384),
    .A1(\cpu.PC[4] ));
 sg13g2_nand3_1 _10083_ (.B(_04387_),
    .C(_04388_),
    .A(_04363_),
    .Y(_04389_));
 sg13g2_mux2_1 _10084_ (.A0(net3003),
    .A1(\cpu.regs[13][4] ),
    .S(net3220),
    .X(_00699_));
 sg13g2_nor2_1 _10085_ (.A(net3261),
    .B(_04133_),
    .Y(_04390_));
 sg13g2_nor2_1 _10086_ (.A(_04240_),
    .B(_04390_),
    .Y(_04391_));
 sg13g2_inv_1 _10087_ (.Y(_04392_),
    .A(_04391_));
 sg13g2_a21oi_1 _10088_ (.A1(net3286),
    .A2(_04392_),
    .Y(_04393_),
    .B1(_04238_));
 sg13g2_mux2_1 _10089_ (.A0(_04277_),
    .A1(_04393_),
    .S(net3278),
    .X(_04394_));
 sg13g2_nand2_1 _10090_ (.Y(_04395_),
    .A(net3305),
    .B(_04394_));
 sg13g2_o21ai_1 _10091_ (.B1(_04395_),
    .Y(_04396_),
    .A1(net3305),
    .A2(_04341_));
 sg13g2_mux2_2 _10092_ (.A0(_04377_),
    .A1(_04396_),
    .S(net3295),
    .X(_04397_));
 sg13g2_nand2_1 _10093_ (.Y(_04398_),
    .A(_03729_),
    .B(_03732_));
 sg13g2_a21o_1 _10094_ (.A2(_04398_),
    .A1(net3375),
    .B1(net3411),
    .X(_04399_));
 sg13g2_o21ai_1 _10095_ (.B1(_04399_),
    .Y(_04400_),
    .A1(_03729_),
    .A2(_03732_));
 sg13g2_o21ai_1 _10096_ (.B1(_04400_),
    .Y(_04401_),
    .A1(net3454),
    .A2(_04398_));
 sg13g2_a21oi_1 _10097_ (.A1(net3353),
    .A2(_04397_),
    .Y(_04402_),
    .B1(_04401_));
 sg13g2_nand2_1 _10098_ (.Y(_04403_),
    .A(net3303),
    .B(_04333_));
 sg13g2_a21oi_1 _10099_ (.A1(net3268),
    .A2(_04170_),
    .Y(_04404_),
    .B1(_04240_));
 sg13g2_nand2_1 _10100_ (.Y(_04405_),
    .A(net3283),
    .B(_04404_));
 sg13g2_o21ai_1 _10101_ (.B1(_04405_),
    .Y(_04406_),
    .A1(net3283),
    .A2(_04176_));
 sg13g2_or2_1 _10102_ (.X(_04407_),
    .B(_04269_),
    .A(net3272));
 sg13g2_o21ai_1 _10103_ (.B1(_04407_),
    .Y(_04408_),
    .A1(net3277),
    .A2(_04406_));
 sg13g2_o21ai_1 _10104_ (.B1(_04403_),
    .Y(_04409_),
    .A1(net3303),
    .A2(_04408_));
 sg13g2_nor2_1 _10105_ (.A(net3290),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_a21oi_2 _10106_ (.B1(_04410_),
    .Y(_04411_),
    .A2(_04368_),
    .A1(net3290));
 sg13g2_a22oi_1 _10107_ (.Y(_04412_),
    .B1(_04411_),
    .B2(net3313),
    .A2(net3338),
    .A1(_04021_));
 sg13g2_a21oi_2 _10108_ (.B1(net3357),
    .Y(_04413_),
    .A2(_04412_),
    .A1(_04402_));
 sg13g2_a221oi_1 _10109_ (.B2(\cpu.PCreg0[5] ),
    .C1(_04413_),
    .B1(net3317),
    .A1(\cpu.PC[5] ),
    .Y(_04414_),
    .A2(net3383));
 sg13g2_nor2_1 _10110_ (.A(net3134),
    .B(net3235),
    .Y(_04415_));
 sg13g2_a22oi_1 _10111_ (.Y(_04416_),
    .B1(_03529_),
    .B2(_04415_),
    .A2(_03525_),
    .A1(net3133));
 sg13g2_nor2_1 _10112_ (.A(net3137),
    .B(_03596_),
    .Y(_04417_));
 sg13g2_a21oi_1 _10113_ (.A1(net3137),
    .A2(\cdi[29] ),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_nor2_1 _10114_ (.A(_02515_),
    .B(_03525_),
    .Y(_04419_));
 sg13g2_a21oi_1 _10115_ (.A1(_02515_),
    .A2(\cdi[21] ),
    .Y(_04420_),
    .B1(_04419_));
 sg13g2_a221oi_1 _10116_ (.B2(_02510_),
    .C1(_01764_),
    .B1(_04420_),
    .A1(_02511_),
    .Y(_04421_),
    .A2(_04418_));
 sg13g2_o21ai_1 _10117_ (.B1(_04421_),
    .Y(_04422_),
    .A1(_02510_),
    .A2(_04416_));
 sg13g2_nand2_2 _10118_ (.Y(_04423_),
    .A(_04414_),
    .B(_04422_));
 sg13g2_mux2_1 _10119_ (.A0(net3030),
    .A1(\cpu.regs[13][5] ),
    .S(net3223),
    .X(_00700_));
 sg13g2_nand2_1 _10120_ (.Y(_04424_),
    .A(_04018_),
    .B(net3338));
 sg13g2_nor2_1 _10121_ (.A(net3305),
    .B(_04375_),
    .Y(_04425_));
 sg13g2_o21ai_1 _10122_ (.B1(net3129),
    .Y(_04426_),
    .A1(net3262),
    .A2(_04187_));
 sg13g2_a21oi_1 _10123_ (.A1(net3285),
    .A2(_04426_),
    .Y(_04427_),
    .B1(_04238_));
 sg13g2_nand2b_1 _10124_ (.Y(_04428_),
    .B(net3275),
    .A_N(_04427_));
 sg13g2_o21ai_1 _10125_ (.B1(_04428_),
    .Y(_04429_),
    .A1(net3275),
    .A2(_04305_));
 sg13g2_a21oi_1 _10126_ (.A1(net3305),
    .A2(_04429_),
    .Y(_04430_),
    .B1(_04425_));
 sg13g2_mux2_2 _10127_ (.A0(_04396_),
    .A1(_04430_),
    .S(net3295),
    .X(_04431_));
 sg13g2_o21ai_1 _10128_ (.B1(net3129),
    .Y(_04432_),
    .A1(net3261),
    .A2(_04194_));
 sg13g2_nor2_1 _10129_ (.A(net3281),
    .B(_04200_),
    .Y(_04433_));
 sg13g2_a21oi_1 _10130_ (.A1(net3281),
    .A2(_04432_),
    .Y(_04434_),
    .B1(_04433_));
 sg13g2_nand2_1 _10131_ (.Y(_04435_),
    .A(net3270),
    .B(_04434_));
 sg13g2_o21ai_1 _10132_ (.B1(_04435_),
    .Y(_04436_),
    .A1(net3270),
    .A2(_04311_));
 sg13g2_nor2_1 _10133_ (.A(net3302),
    .B(_04436_),
    .Y(_04437_));
 sg13g2_a21oi_1 _10134_ (.A1(net3302),
    .A2(_04367_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_nor2b_1 _10135_ (.A(net3290),
    .B_N(_04438_),
    .Y(_04439_));
 sg13g2_a21oi_2 _10136_ (.B1(_04439_),
    .Y(_04440_),
    .A2(_04409_),
    .A1(net3289));
 sg13g2_nor2_1 _10137_ (.A(_03718_),
    .B(_03721_),
    .Y(_04441_));
 sg13g2_nand2_1 _10138_ (.Y(_04442_),
    .A(_03718_),
    .B(_03721_));
 sg13g2_a21oi_1 _10139_ (.A1(net3374),
    .A2(_04442_),
    .Y(_04443_),
    .B1(net3411));
 sg13g2_nor2_1 _10140_ (.A(net3454),
    .B(_04442_),
    .Y(_04444_));
 sg13g2_o21ai_1 _10141_ (.B1(_04424_),
    .Y(_04445_),
    .A1(net3311),
    .A2(_04440_));
 sg13g2_a21oi_1 _10142_ (.A1(net3352),
    .A2(_04431_),
    .Y(_04446_),
    .B1(_04444_));
 sg13g2_o21ai_1 _10143_ (.B1(_04446_),
    .Y(_04447_),
    .A1(_04441_),
    .A2(_04443_));
 sg13g2_o21ai_1 _10144_ (.B1(net3356),
    .Y(_04448_),
    .A1(_04445_),
    .A2(_04447_));
 sg13g2_a22oi_1 _10145_ (.Y(_04449_),
    .B1(net3317),
    .B2(\cpu.PCreg0[6] ),
    .A2(net3384),
    .A1(\cpu.PC[6] ));
 sg13g2_a21oi_1 _10146_ (.A1(net3137),
    .A2(\cdi[30] ),
    .Y(_04450_),
    .B1(_02512_));
 sg13g2_o21ai_1 _10147_ (.B1(_04450_),
    .Y(_04451_),
    .A1(net3137),
    .A2(_03605_));
 sg13g2_nand3_1 _10148_ (.B(_03542_),
    .C(_04260_),
    .A(_03539_),
    .Y(_04452_));
 sg13g2_or2_1 _10149_ (.X(_04453_),
    .B(\cdi[6] ),
    .A(_02518_));
 sg13g2_nand4_1 _10150_ (.B(_04451_),
    .C(_04452_),
    .A(net3448),
    .Y(_04454_),
    .D(_04453_));
 sg13g2_nand3_1 _10151_ (.B(_04449_),
    .C(_04454_),
    .A(_04448_),
    .Y(_04455_));
 sg13g2_mux2_1 _10152_ (.A0(net3038),
    .A1(\cpu.regs[13][6] ),
    .S(net3220),
    .X(_00701_));
 sg13g2_nor3_1 _10153_ (.A(net3137),
    .B(net3235),
    .C(\cdi[7] ),
    .Y(_04456_));
 sg13g2_nor2b_1 _10154_ (.A(\cdi[23] ),
    .B_N(_04415_),
    .Y(_04457_));
 sg13g2_o21ai_1 _10155_ (.B1(net3459),
    .Y(_04458_),
    .A1(_04456_),
    .A2(_04457_));
 sg13g2_mux2_1 _10156_ (.A0(_03609_),
    .A1(_03611_),
    .S(net3137),
    .X(_04459_));
 sg13g2_nand2_1 _10157_ (.Y(_04460_),
    .A(_02511_),
    .B(_04459_));
 sg13g2_nand2_1 _10158_ (.Y(_04461_),
    .A(_04458_),
    .B(_04460_));
 sg13g2_mux2_1 _10159_ (.A0(\cdi[7] ),
    .A1(\cdi[23] ),
    .S(_02515_),
    .X(_04462_));
 sg13g2_o21ai_1 _10160_ (.B1(net3448),
    .Y(_04463_),
    .A1(net3459),
    .A2(_04462_));
 sg13g2_nand2_1 _10161_ (.Y(_04464_),
    .A(net3276),
    .B(_04331_));
 sg13g2_o21ai_1 _10162_ (.B1(net3129),
    .Y(_04465_),
    .A1(net3262),
    .A2(_04143_));
 sg13g2_nor2_1 _10163_ (.A(net3285),
    .B(_04465_),
    .Y(_04466_));
 sg13g2_a21oi_1 _10164_ (.A1(net3285),
    .A2(_04152_),
    .Y(_04467_),
    .B1(_04466_));
 sg13g2_o21ai_1 _10165_ (.B1(_04464_),
    .Y(_04468_),
    .A1(net3276),
    .A2(_04467_));
 sg13g2_nand2_1 _10166_ (.Y(_04469_),
    .A(net3305),
    .B(_04408_));
 sg13g2_o21ai_1 _10167_ (.B1(_04469_),
    .Y(_04470_),
    .A1(net3301),
    .A2(_04468_));
 sg13g2_nand2_1 _10168_ (.Y(_04471_),
    .A(net3290),
    .B(_04438_));
 sg13g2_o21ai_1 _10169_ (.B1(_04471_),
    .Y(_04472_),
    .A1(net3290),
    .A2(_04470_));
 sg13g2_a21oi_1 _10170_ (.A1(net3269),
    .A2(_04158_),
    .Y(_04473_),
    .B1(_04240_));
 sg13g2_o21ai_1 _10171_ (.B1(_04239_),
    .Y(_04474_),
    .A1(net3282),
    .A2(_04473_));
 sg13g2_nand2_1 _10172_ (.Y(_04475_),
    .A(net3272),
    .B(_04340_));
 sg13g2_o21ai_1 _10173_ (.B1(_04475_),
    .Y(_04476_),
    .A1(net3270),
    .A2(_04474_));
 sg13g2_mux2_1 _10174_ (.A0(_04394_),
    .A1(_04476_),
    .S(net3305),
    .X(_04477_));
 sg13g2_mux2_1 _10175_ (.A0(_04430_),
    .A1(_04477_),
    .S(net3295),
    .X(_04478_));
 sg13g2_nand2_1 _10176_ (.Y(_04479_),
    .A(_03707_),
    .B(_03710_));
 sg13g2_a21o_1 _10177_ (.A2(_04479_),
    .A1(net3374),
    .B1(net3411),
    .X(_04480_));
 sg13g2_o21ai_1 _10178_ (.B1(_04480_),
    .Y(_04481_),
    .A1(_03707_),
    .A2(_03710_));
 sg13g2_o21ai_1 _10179_ (.B1(_04481_),
    .Y(_04482_),
    .A1(net3454),
    .A2(_04479_));
 sg13g2_a221oi_1 _10180_ (.B2(net3352),
    .C1(_04482_),
    .B1(_04478_),
    .A1(net3313),
    .Y(_04483_),
    .A2(_04472_));
 sg13g2_o21ai_1 _10181_ (.B1(_04483_),
    .Y(_04484_),
    .A1(_04037_),
    .A2(net3378));
 sg13g2_and2_1 _10182_ (.A(\cpu.PC[7] ),
    .B(net3383),
    .X(_04485_));
 sg13g2_a221oi_1 _10183_ (.B2(_04115_),
    .C1(_04485_),
    .B1(_04484_),
    .A1(\cpu.PCreg0[7] ),
    .Y(_04486_),
    .A2(net3317));
 sg13g2_o21ai_1 _10184_ (.B1(_04486_),
    .Y(_04487_),
    .A1(_04461_),
    .A2(_04463_));
 sg13g2_mux2_1 _10185_ (.A0(net3045),
    .A1(\cpu.regs[13][7] ),
    .S(net3222),
    .X(_00702_));
 sg13g2_nand3b_1 _10186_ (.B(_04458_),
    .C(_04460_),
    .Y(_04488_),
    .A_N(net3694));
 sg13g2_a21oi_1 _10187_ (.A1(net3459),
    .A2(_04488_),
    .Y(_04489_),
    .B1(_01764_));
 sg13g2_a21oi_1 _10188_ (.A1(_02506_),
    .A2(\cdi[24] ),
    .Y(_04490_),
    .B1(net3459));
 sg13g2_o21ai_1 _10189_ (.B1(_04490_),
    .Y(_04491_),
    .A1(_02506_),
    .A2(_03567_));
 sg13g2_nand2_1 _10190_ (.Y(_04492_),
    .A(net3043),
    .B(_04491_));
 sg13g2_nor2_1 _10191_ (.A(net3275),
    .B(_04373_),
    .Y(_04493_));
 sg13g2_o21ai_1 _10192_ (.B1(_04241_),
    .Y(_04494_),
    .A1(net3266),
    .A2(_04216_));
 sg13g2_nor2_1 _10193_ (.A(net3282),
    .B(_04494_),
    .Y(_04495_));
 sg13g2_a21oi_1 _10194_ (.A1(net3282),
    .A2(_04242_),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_a21oi_1 _10195_ (.A1(net3275),
    .A2(_04496_),
    .Y(_04497_),
    .B1(_04493_));
 sg13g2_nand2_1 _10196_ (.Y(_04498_),
    .A(net3301),
    .B(_04497_));
 sg13g2_o21ai_1 _10197_ (.B1(_04498_),
    .Y(_04499_),
    .A1(net3301),
    .A2(_04429_));
 sg13g2_mux2_2 _10198_ (.A0(_04477_),
    .A1(_04499_),
    .S(net3293),
    .X(_04500_));
 sg13g2_nand2_1 _10199_ (.Y(_04501_),
    .A(_03812_),
    .B(_03814_));
 sg13g2_a21o_1 _10200_ (.A2(_04501_),
    .A1(net3374),
    .B1(net3411),
    .X(_04502_));
 sg13g2_o21ai_1 _10201_ (.B1(_04502_),
    .Y(_04503_),
    .A1(_03812_),
    .A2(_03814_));
 sg13g2_o21ai_1 _10202_ (.B1(_04503_),
    .Y(_04504_),
    .A1(net3454),
    .A2(_04501_));
 sg13g2_mux2_1 _10203_ (.A0(_04224_),
    .A1(_04494_),
    .S(net3283),
    .X(_04505_));
 sg13g2_mux2_1 _10204_ (.A0(_04365_),
    .A1(_04505_),
    .S(net3270),
    .X(_04506_));
 sg13g2_nand2_1 _10205_ (.Y(_04507_),
    .A(net3302),
    .B(_04436_));
 sg13g2_o21ai_1 _10206_ (.B1(_04507_),
    .Y(_04508_),
    .A1(net3302),
    .A2(_04506_));
 sg13g2_nand2_1 _10207_ (.Y(_04509_),
    .A(net3294),
    .B(_04470_));
 sg13g2_o21ai_1 _10208_ (.B1(_04509_),
    .Y(_04510_),
    .A1(net3290),
    .A2(_04508_));
 sg13g2_a221oi_1 _10209_ (.B2(net3353),
    .C1(_04504_),
    .B1(_04500_),
    .A1(_04019_),
    .Y(_04511_),
    .A2(net3337));
 sg13g2_o21ai_1 _10210_ (.B1(_04511_),
    .Y(_04512_),
    .A1(net3311),
    .A2(_04510_));
 sg13g2_nand2_1 _10211_ (.Y(_04513_),
    .A(net3356),
    .B(_04512_));
 sg13g2_a22oi_1 _10212_ (.Y(_04514_),
    .B1(net3317),
    .B2(\cpu.PCreg0[8] ),
    .A2(net3383),
    .A1(\cpu.PC[8] ));
 sg13g2_nand3_1 _10213_ (.B(_04513_),
    .C(_04514_),
    .A(_04492_),
    .Y(_04515_));
 sg13g2_mux2_1 _10214_ (.A0(net3028),
    .A1(\cpu.regs[13][8] ),
    .S(net3222),
    .X(_00703_));
 sg13g2_nor2_1 _10215_ (.A(_04030_),
    .B(net3378),
    .Y(_04516_));
 sg13g2_nand2b_1 _10216_ (.Y(_04517_),
    .B(net3281),
    .A_N(_04276_));
 sg13g2_o21ai_1 _10217_ (.B1(_04517_),
    .Y(_04518_),
    .A1(net3281),
    .A2(_04465_));
 sg13g2_mux2_1 _10218_ (.A0(_04393_),
    .A1(_04518_),
    .S(net3274),
    .X(_04519_));
 sg13g2_nor2b_1 _10219_ (.A(net3301),
    .B_N(_04476_),
    .Y(_04520_));
 sg13g2_a21oi_2 _10220_ (.B1(_04520_),
    .Y(_04521_),
    .A2(_04519_),
    .A1(net3302));
 sg13g2_nor2_1 _10221_ (.A(net3293),
    .B(_04499_),
    .Y(_04522_));
 sg13g2_a21oi_2 _10222_ (.B1(_04522_),
    .Y(_04523_),
    .A2(_04521_),
    .A1(net3293));
 sg13g2_nand2_1 _10223_ (.Y(_04524_),
    .A(net3348),
    .B(_04523_));
 sg13g2_nor2_1 _10224_ (.A(net3284),
    .B(_04268_),
    .Y(_04525_));
 sg13g2_a21oi_1 _10225_ (.A1(net3282),
    .A2(_04473_),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_nor2_1 _10226_ (.A(net3271),
    .B(_04406_),
    .Y(_04527_));
 sg13g2_a21oi_1 _10227_ (.A1(net3271),
    .A2(_04526_),
    .Y(_04528_),
    .B1(_04527_));
 sg13g2_nor2b_1 _10228_ (.A(net3298),
    .B_N(_04528_),
    .Y(_04529_));
 sg13g2_a21oi_1 _10229_ (.A1(net3301),
    .A2(_04468_),
    .Y(_04530_),
    .B1(_04529_));
 sg13g2_nor2_1 _10230_ (.A(net3294),
    .B(_04530_),
    .Y(_04531_));
 sg13g2_a21oi_2 _10231_ (.B1(_04531_),
    .Y(_04532_),
    .A2(_04508_),
    .A1(net3294));
 sg13g2_nor2_1 _10232_ (.A(net3310),
    .B(_04532_),
    .Y(_04533_));
 sg13g2_or2_1 _10233_ (.X(_04534_),
    .B(_03822_),
    .A(_03819_));
 sg13g2_nand2_1 _10234_ (.Y(_04535_),
    .A(net3374),
    .B(_04534_));
 sg13g2_a22oi_1 _10235_ (.Y(_04536_),
    .B1(net3409),
    .B2(_04535_),
    .A2(_03822_),
    .A1(_03819_));
 sg13g2_o21ai_1 _10236_ (.B1(_04524_),
    .Y(_04537_),
    .A1(net3454),
    .A2(_04534_));
 sg13g2_nor4_1 _10237_ (.A(_04516_),
    .B(_04533_),
    .C(_04536_),
    .D(_04537_),
    .Y(_04538_));
 sg13g2_nor2_1 _10238_ (.A(net3357),
    .B(_04538_),
    .Y(_04539_));
 sg13g2_a221oi_1 _10239_ (.B2(\cpu.PCreg0[9] ),
    .C1(_04539_),
    .B1(net3318),
    .A1(\cpu.PC[9] ),
    .Y(_04540_),
    .A2(net3383));
 sg13g2_nor2_1 _10240_ (.A(_02514_),
    .B(_04294_),
    .Y(_04541_));
 sg13g2_o21ai_1 _10241_ (.B1(net3043),
    .Y(_04542_),
    .A1(net3624),
    .A2(\cdi[9] ));
 sg13g2_o21ai_1 _10242_ (.B1(_04540_),
    .Y(_04543_),
    .A1(_04541_),
    .A2(_04542_));
 sg13g2_mux2_1 _10243_ (.A0(net3026),
    .A1(\cpu.regs[13][9] ),
    .S(net3222),
    .X(_00704_));
 sg13g2_nor2_1 _10244_ (.A(_04035_),
    .B(net3378),
    .Y(_04544_));
 sg13g2_nor2_1 _10245_ (.A(net3282),
    .B(_04432_),
    .Y(_04545_));
 sg13g2_a21oi_1 _10246_ (.A1(net3281),
    .A2(_04303_),
    .Y(_04546_),
    .B1(_04545_));
 sg13g2_nand2_1 _10247_ (.Y(_04547_),
    .A(net3274),
    .B(_04546_));
 sg13g2_o21ai_1 _10248_ (.B1(_04547_),
    .Y(_04548_),
    .A1(net3274),
    .A2(_04427_));
 sg13g2_nand2_1 _10249_ (.Y(_04549_),
    .A(net3300),
    .B(_04548_));
 sg13g2_o21ai_1 _10250_ (.B1(_04549_),
    .Y(_04550_),
    .A1(net3301),
    .A2(_04497_));
 sg13g2_nand2b_1 _10251_ (.Y(_04551_),
    .B(net3291),
    .A_N(_04550_));
 sg13g2_o21ai_1 _10252_ (.B1(_04551_),
    .Y(_04552_),
    .A1(net3292),
    .A2(_04521_));
 sg13g2_and2_1 _10253_ (.A(net3354),
    .B(_04552_),
    .X(_04553_));
 sg13g2_nand2_1 _10254_ (.Y(_04554_),
    .A(net3274),
    .B(_04434_));
 sg13g2_nand2_1 _10255_ (.Y(_04555_),
    .A(net3281),
    .B(_04426_));
 sg13g2_o21ai_1 _10256_ (.B1(_04555_),
    .Y(_04556_),
    .A1(net3282),
    .A2(_04309_));
 sg13g2_o21ai_1 _10257_ (.B1(_04554_),
    .Y(_04557_),
    .A1(net3274),
    .A2(_04556_));
 sg13g2_nand2_1 _10258_ (.Y(_04558_),
    .A(net3298),
    .B(_04506_));
 sg13g2_o21ai_1 _10259_ (.B1(_04558_),
    .Y(_04559_),
    .A1(net3298),
    .A2(_04557_));
 sg13g2_nor2b_1 _10260_ (.A(net3294),
    .B_N(_04559_),
    .Y(_04560_));
 sg13g2_a21oi_2 _10261_ (.B1(_04560_),
    .Y(_04561_),
    .A2(_04530_),
    .A1(net3294));
 sg13g2_nand2_1 _10262_ (.Y(_04562_),
    .A(net3313),
    .B(_04561_));
 sg13g2_nand2b_1 _10263_ (.Y(_04563_),
    .B(_03796_),
    .A_N(_03794_));
 sg13g2_nand2_1 _10264_ (.Y(_04564_),
    .A(net3373),
    .B(_04563_));
 sg13g2_a22oi_1 _10265_ (.Y(_04565_),
    .B1(net3408),
    .B2(_04564_),
    .A2(_03797_),
    .A1(_03794_));
 sg13g2_o21ai_1 _10266_ (.B1(_04562_),
    .Y(_04566_),
    .A1(net3452),
    .A2(_04563_));
 sg13g2_nor4_2 _10267_ (.A(_04544_),
    .B(_04553_),
    .C(_04565_),
    .Y(_04567_),
    .D(_04566_));
 sg13g2_nor2_1 _10268_ (.A(net3358),
    .B(_04567_),
    .Y(_04568_));
 sg13g2_a221oi_1 _10269_ (.B2(\cpu.PCreg0[10] ),
    .C1(_04568_),
    .B1(net3317),
    .A1(\cpu.PC[10] ),
    .Y(_04569_),
    .A2(net3383));
 sg13g2_nor2_1 _10270_ (.A(_02514_),
    .B(_04299_),
    .Y(_04570_));
 sg13g2_o21ai_1 _10271_ (.B1(net3043),
    .Y(_04571_),
    .A1(net3625),
    .A2(\cdi[10] ));
 sg13g2_o21ai_1 _10272_ (.B1(_04569_),
    .Y(_04572_),
    .A1(_04570_),
    .A2(_04571_));
 sg13g2_mux2_1 _10273_ (.A0(net3024),
    .A1(\cpu.regs[13][10] ),
    .S(net3223),
    .X(_00705_));
 sg13g2_a22oi_1 _10274_ (.Y(_04573_),
    .B1(_04328_),
    .B2(_02513_),
    .A2(_03588_),
    .A1(net3695));
 sg13g2_nor2_1 _10275_ (.A(net3286),
    .B(_04339_),
    .Y(_04574_));
 sg13g2_a21oi_1 _10276_ (.A1(net3285),
    .A2(_04404_),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_mux2_1 _10277_ (.A0(_04474_),
    .A1(_04575_),
    .S(net3278),
    .X(_04576_));
 sg13g2_nand2_1 _10278_ (.Y(_04577_),
    .A(net3300),
    .B(_04576_));
 sg13g2_o21ai_1 _10279_ (.B1(_04577_),
    .Y(_04578_),
    .A1(net3300),
    .A2(_04519_));
 sg13g2_nor2b_1 _10280_ (.A(net3291),
    .B_N(_04550_),
    .Y(_04579_));
 sg13g2_a21oi_2 _10281_ (.B1(_04579_),
    .Y(_04580_),
    .A2(_04578_),
    .A1(net3291));
 sg13g2_nor2_1 _10282_ (.A(net3285),
    .B(_04391_),
    .Y(_04581_));
 sg13g2_a21oi_1 _10283_ (.A1(net3285),
    .A2(_04329_),
    .Y(_04582_),
    .B1(_04581_));
 sg13g2_nor2_1 _10284_ (.A(net3274),
    .B(_04582_),
    .Y(_04583_));
 sg13g2_a21oi_1 _10285_ (.A1(net3274),
    .A2(_04467_),
    .Y(_04584_),
    .B1(_04583_));
 sg13g2_nand2b_1 _10286_ (.Y(_04585_),
    .B(net3298),
    .A_N(_04528_));
 sg13g2_o21ai_1 _10287_ (.B1(_04585_),
    .Y(_04586_),
    .A1(net3298),
    .A2(_04584_));
 sg13g2_mux2_1 _10288_ (.A0(_04586_),
    .A1(_04559_),
    .S(net3294),
    .X(_04587_));
 sg13g2_or2_1 _10289_ (.X(_04588_),
    .B(_03804_),
    .A(_03803_));
 sg13g2_nand2_1 _10290_ (.Y(_04589_),
    .A(_03803_),
    .B(_03804_));
 sg13g2_a21o_1 _10291_ (.A2(_04589_),
    .A1(net3372),
    .B1(net3410),
    .X(_04590_));
 sg13g2_nor2_1 _10292_ (.A(net3452),
    .B(_04589_),
    .Y(_04591_));
 sg13g2_a21oi_1 _10293_ (.A1(_04588_),
    .A2(_04590_),
    .Y(_04592_),
    .B1(_04591_));
 sg13g2_o21ai_1 _10294_ (.B1(_04592_),
    .Y(_04593_),
    .A1(net3310),
    .A2(_04587_));
 sg13g2_a221oi_1 _10295_ (.B2(net3348),
    .C1(_04593_),
    .B1(_04580_),
    .A1(_04001_),
    .Y(_04594_),
    .A2(net3337));
 sg13g2_a22oi_1 _10296_ (.Y(_04595_),
    .B1(net3314),
    .B2(\cpu.PCreg0[11] ),
    .A2(net3381),
    .A1(\cpu.PC[11] ));
 sg13g2_o21ai_1 _10297_ (.B1(_04595_),
    .Y(_04596_),
    .A1(net3358),
    .A2(_04594_));
 sg13g2_a21o_2 _10298_ (.A2(_04573_),
    .A1(_04489_),
    .B1(_04596_),
    .X(_04597_));
 sg13g2_mux2_1 _10299_ (.A0(net3022),
    .A1(\cpu.regs[13][11] ),
    .S(net3223),
    .X(_00706_));
 sg13g2_nand2_1 _10300_ (.Y(_04598_),
    .A(_02515_),
    .B(\cdi[28] ));
 sg13g2_o21ai_1 _10301_ (.B1(_04598_),
    .Y(_04599_),
    .A1(_02506_),
    .A2(_03593_));
 sg13g2_o21ai_1 _10302_ (.B1(net3043),
    .Y(_04600_),
    .A1(net3459),
    .A2(_04599_));
 sg13g2_mux2_1 _10303_ (.A0(_04364_),
    .A1(_04372_),
    .S(net3282),
    .X(_04601_));
 sg13g2_mux2_1 _10304_ (.A0(_04496_),
    .A1(_04601_),
    .S(net3275),
    .X(_04602_));
 sg13g2_mux2_1 _10305_ (.A0(_04548_),
    .A1(_04602_),
    .S(net3299),
    .X(_04603_));
 sg13g2_nand2b_1 _10306_ (.Y(_04604_),
    .B(net3291),
    .A_N(_04603_));
 sg13g2_o21ai_1 _10307_ (.B1(_04604_),
    .Y(_04605_),
    .A1(net3291),
    .A2(_04578_));
 sg13g2_mux2_1 _10308_ (.A0(_04505_),
    .A1(_04601_),
    .S(net3270),
    .X(_04606_));
 sg13g2_nor2_1 _10309_ (.A(net3298),
    .B(_04606_),
    .Y(_04607_));
 sg13g2_a21oi_1 _10310_ (.A1(net3298),
    .A2(_04557_),
    .Y(_04608_),
    .B1(_04607_));
 sg13g2_mux2_1 _10311_ (.A0(_04608_),
    .A1(_04586_),
    .S(net3294),
    .X(_04609_));
 sg13g2_nand2b_1 _10312_ (.Y(_04610_),
    .B(_03788_),
    .A_N(_03786_));
 sg13g2_nand2_1 _10313_ (.Y(_04611_),
    .A(net3373),
    .B(_04610_));
 sg13g2_a22oi_1 _10314_ (.Y(_04612_),
    .B1(net3408),
    .B2(_04611_),
    .A2(_03789_),
    .A1(_03786_));
 sg13g2_nor2_1 _10315_ (.A(net3452),
    .B(_04610_),
    .Y(_04613_));
 sg13g2_nor2_1 _10316_ (.A(_04612_),
    .B(_04613_),
    .Y(_04614_));
 sg13g2_o21ai_1 _10317_ (.B1(_04614_),
    .Y(_04615_),
    .A1(net3310),
    .A2(_04609_));
 sg13g2_a221oi_1 _10318_ (.B2(net3348),
    .C1(_04615_),
    .B1(_04605_),
    .A1(_04044_),
    .Y(_04616_),
    .A2(net3337));
 sg13g2_a22oi_1 _10319_ (.Y(_04617_),
    .B1(net3314),
    .B2(\cpu.PCreg0[12] ),
    .A2(net3381),
    .A1(\cpu.PC[12] ));
 sg13g2_o21ai_1 _10320_ (.B1(_04617_),
    .Y(_04618_),
    .A1(net3358),
    .A2(_04616_));
 sg13g2_nand2b_1 _10321_ (.Y(_04619_),
    .B(_04600_),
    .A_N(_04618_));
 sg13g2_mux2_1 _10322_ (.A0(net3001),
    .A1(\cpu.regs[13][12] ),
    .S(net3220),
    .X(_00707_));
 sg13g2_a22oi_1 _10323_ (.Y(_04620_),
    .B1(_04418_),
    .B2(_02513_),
    .A2(_03596_),
    .A1(net3698));
 sg13g2_nand2_2 _10324_ (.Y(_04621_),
    .A(net3043),
    .B(_04620_));
 sg13g2_mux2_1 _10325_ (.A0(_04518_),
    .A1(_04582_),
    .S(net3275),
    .X(_04622_));
 sg13g2_nor2_1 _10326_ (.A(net3300),
    .B(_04576_),
    .Y(_04623_));
 sg13g2_a21oi_2 _10327_ (.B1(_04623_),
    .Y(_04624_),
    .A2(_04622_),
    .A1(net3300));
 sg13g2_nor2b_1 _10328_ (.A(net3291),
    .B_N(_04603_),
    .Y(_04625_));
 sg13g2_a21oi_2 _10329_ (.B1(_04625_),
    .Y(_04626_),
    .A2(_04624_),
    .A1(net3291));
 sg13g2_mux2_1 _10330_ (.A0(_04526_),
    .A1(_04575_),
    .S(net3271),
    .X(_04627_));
 sg13g2_nor2_1 _10331_ (.A(net3299),
    .B(_04627_),
    .Y(_04628_));
 sg13g2_a21oi_1 _10332_ (.A1(net3298),
    .A2(_04584_),
    .Y(_04629_),
    .B1(_04628_));
 sg13g2_mux2_1 _10333_ (.A0(_04629_),
    .A1(_04608_),
    .S(net3294),
    .X(_04630_));
 sg13g2_nor2_1 _10334_ (.A(net3310),
    .B(_04630_),
    .Y(_04631_));
 sg13g2_nand2b_1 _10335_ (.Y(_04632_),
    .B(_03780_),
    .A_N(_03778_));
 sg13g2_inv_1 _10336_ (.Y(_04633_),
    .A(_04632_));
 sg13g2_nand2_1 _10337_ (.Y(_04634_),
    .A(net3373),
    .B(_04632_));
 sg13g2_a22oi_1 _10338_ (.Y(_04635_),
    .B1(net3408),
    .B2(_04634_),
    .A2(_03781_),
    .A1(_03778_));
 sg13g2_a221oi_1 _10339_ (.B2(_04253_),
    .C1(_04635_),
    .B1(_04633_),
    .A1(net3348),
    .Y(_04636_),
    .A2(_04626_));
 sg13g2_o21ai_1 _10340_ (.B1(_04636_),
    .Y(_04637_),
    .A1(_04051_),
    .A2(net3377));
 sg13g2_o21ai_1 _10341_ (.B1(net3356),
    .Y(_04638_),
    .A1(_04631_),
    .A2(_04637_));
 sg13g2_a22oi_1 _10342_ (.Y(_04639_),
    .B1(net3314),
    .B2(\cpu.PCreg0[13] ),
    .A2(net3381),
    .A1(\cpu.PC[13] ));
 sg13g2_nand3_1 _10343_ (.B(_04638_),
    .C(_04639_),
    .A(_04621_),
    .Y(_04640_));
 sg13g2_mux2_1 _10344_ (.A0(net3020),
    .A1(\cpu.regs[13][13] ),
    .S(net3220),
    .X(_00708_));
 sg13g2_a21oi_1 _10345_ (.A1(_02515_),
    .A2(\cdi[30] ),
    .Y(_04641_),
    .B1(net3459));
 sg13g2_o21ai_1 _10346_ (.B1(_04641_),
    .Y(_04642_),
    .A1(_02506_),
    .A2(_03605_));
 sg13g2_or2_1 _10347_ (.X(_04643_),
    .B(_04556_),
    .A(net3271));
 sg13g2_o21ai_1 _10348_ (.B1(_04643_),
    .Y(_04644_),
    .A1(net3274),
    .A2(_04546_));
 sg13g2_nor2_1 _10349_ (.A(net3299),
    .B(_04602_),
    .Y(_04645_));
 sg13g2_a21oi_1 _10350_ (.A1(net3299),
    .A2(_04644_),
    .Y(_04646_),
    .B1(_04645_));
 sg13g2_mux2_1 _10351_ (.A0(_04624_),
    .A1(_04646_),
    .S(net3291),
    .X(_04647_));
 sg13g2_nor2_1 _10352_ (.A(net3299),
    .B(_04644_),
    .Y(_04648_));
 sg13g2_a21oi_1 _10353_ (.A1(net3299),
    .A2(_04606_),
    .Y(_04649_),
    .B1(_04648_));
 sg13g2_nand2_1 _10354_ (.Y(_04650_),
    .A(net3292),
    .B(_04629_));
 sg13g2_o21ai_1 _10355_ (.B1(_04650_),
    .Y(_04651_),
    .A1(net3292),
    .A2(_04649_));
 sg13g2_nor2_1 _10356_ (.A(net3310),
    .B(_04651_),
    .Y(_04652_));
 sg13g2_nand2_1 _10357_ (.Y(_04653_),
    .A(_03762_),
    .B(_03764_));
 sg13g2_a21o_1 _10358_ (.A2(_04653_),
    .A1(net3372),
    .B1(net3410),
    .X(_04654_));
 sg13g2_o21ai_1 _10359_ (.B1(_04654_),
    .Y(_04655_),
    .A1(_03762_),
    .A2(_03764_));
 sg13g2_o21ai_1 _10360_ (.B1(_04655_),
    .Y(_04656_),
    .A1(net3453),
    .A2(_04653_));
 sg13g2_nor2_1 _10361_ (.A(_04652_),
    .B(_04656_),
    .Y(_04657_));
 sg13g2_o21ai_1 _10362_ (.B1(_04657_),
    .Y(_04658_),
    .A1(net3340),
    .A2(_04647_));
 sg13g2_a21oi_1 _10363_ (.A1(_03991_),
    .A2(net3337),
    .Y(_04659_),
    .B1(_04658_));
 sg13g2_a22oi_1 _10364_ (.Y(_04660_),
    .B1(net3314),
    .B2(\cpu.PCreg0[14] ),
    .A2(net3381),
    .A1(\cpu.PC[14] ));
 sg13g2_o21ai_1 _10365_ (.B1(_04660_),
    .Y(_04661_),
    .A1(net3358),
    .A2(_04659_));
 sg13g2_a21oi_2 _10366_ (.B1(_04661_),
    .Y(_04662_),
    .A2(_04642_),
    .A1(net3043));
 sg13g2_nand2_1 _10367_ (.Y(_04663_),
    .A(\cpu.regs[13][14] ),
    .B(net3222));
 sg13g2_o21ai_1 _10368_ (.B1(_04663_),
    .Y(_00709_),
    .A1(net3222),
    .A2(net3036));
 sg13g2_nor2_1 _10369_ (.A(_03990_),
    .B(net3377),
    .Y(_04664_));
 sg13g2_nor2_1 _10370_ (.A(net3299),
    .B(_04622_),
    .Y(_04665_));
 sg13g2_a21oi_1 _10371_ (.A1(net3299),
    .A2(_04627_),
    .Y(_04666_),
    .B1(_04665_));
 sg13g2_nor2_1 _10372_ (.A(net3292),
    .B(_04646_),
    .Y(_04667_));
 sg13g2_a21oi_1 _10373_ (.A1(net3292),
    .A2(_04666_),
    .Y(_04668_),
    .B1(_04667_));
 sg13g2_nor2_1 _10374_ (.A(net3339),
    .B(_04668_),
    .Y(_04669_));
 sg13g2_nand2b_1 _10375_ (.Y(_04670_),
    .B(_03771_),
    .A_N(_03769_));
 sg13g2_nor2_1 _10376_ (.A(net3453),
    .B(_04670_),
    .Y(_04671_));
 sg13g2_nand2_1 _10377_ (.Y(_04672_),
    .A(net3372),
    .B(_04670_));
 sg13g2_a22oi_1 _10378_ (.Y(_04673_),
    .B1(net3408),
    .B2(_04672_),
    .A2(_03772_),
    .A1(_03769_));
 sg13g2_nor3_1 _10379_ (.A(_04669_),
    .B(_04671_),
    .C(_04673_),
    .Y(_04674_));
 sg13g2_nor2b_1 _10380_ (.A(net3292),
    .B_N(_04666_),
    .Y(_04675_));
 sg13g2_a21oi_1 _10381_ (.A1(net3292),
    .A2(_04649_),
    .Y(_04676_),
    .B1(_04675_));
 sg13g2_o21ai_1 _10382_ (.B1(_04674_),
    .Y(_04677_),
    .A1(net3310),
    .A2(_04676_));
 sg13g2_o21ai_1 _10383_ (.B1(net3355),
    .Y(_04678_),
    .A1(_04664_),
    .A2(_04677_));
 sg13g2_a22oi_1 _10384_ (.Y(_04679_),
    .B1(net3315),
    .B2(\cpu.PCreg0[15] ),
    .A2(net3382),
    .A1(\cpu.PC[15] ));
 sg13g2_nand2_2 _10385_ (.Y(_04680_),
    .A(_04678_),
    .B(_04679_));
 sg13g2_nand2_1 _10386_ (.Y(_04681_),
    .A(_02513_),
    .B(_04459_));
 sg13g2_a22oi_1 _10387_ (.Y(_04682_),
    .B1(_04459_),
    .B2(_02513_),
    .A2(_03609_),
    .A1(net3698));
 sg13g2_a21oi_2 _10388_ (.B1(_04680_),
    .Y(_04683_),
    .A2(_04682_),
    .A1(net3043));
 sg13g2_nand2_1 _10389_ (.Y(_04684_),
    .A(\cpu.regs[13][15] ),
    .B(net3222));
 sg13g2_o21ai_1 _10390_ (.B1(_04684_),
    .Y(_00710_),
    .A1(net3222),
    .A2(net3034));
 sg13g2_nand2_1 _10391_ (.Y(_04685_),
    .A(_02513_),
    .B(_04488_));
 sg13g2_nand3_1 _10392_ (.B(_04681_),
    .C(_04685_),
    .A(net3043),
    .Y(_04686_));
 sg13g2_a21oi_1 _10393_ (.A1(net3695),
    .A2(_03458_),
    .Y(_04687_),
    .B1(net3032));
 sg13g2_nand2_1 _10394_ (.Y(_04688_),
    .A(_04031_),
    .B(net3337));
 sg13g2_nor2_1 _10395_ (.A(net3310),
    .B(_04668_),
    .Y(_04689_));
 sg13g2_nand2_1 _10396_ (.Y(_04690_),
    .A(_03880_),
    .B(_03883_));
 sg13g2_a21o_1 _10397_ (.A2(_04690_),
    .A1(net3371),
    .B1(net3412),
    .X(_04691_));
 sg13g2_o21ai_1 _10398_ (.B1(_04691_),
    .Y(_04692_),
    .A1(_03880_),
    .A2(_03883_));
 sg13g2_o21ai_1 _10399_ (.B1(_04692_),
    .Y(_04693_),
    .A1(net3453),
    .A2(_04690_));
 sg13g2_o21ai_1 _10400_ (.B1(_04688_),
    .Y(_04694_),
    .A1(net3339),
    .A2(_04676_));
 sg13g2_nor3_2 _10401_ (.A(_04689_),
    .B(_04693_),
    .C(_04694_),
    .Y(_04695_));
 sg13g2_a22oi_1 _10402_ (.Y(_04696_),
    .B1(net3314),
    .B2(\cpu.PCreg0[16] ),
    .A2(net3381),
    .A1(\cpu.PC[16] ));
 sg13g2_o21ai_1 _10403_ (.B1(_04696_),
    .Y(_04697_),
    .A1(net3358),
    .A2(_04695_));
 sg13g2_or2_1 _10404_ (.X(_04698_),
    .B(_04697_),
    .A(_04687_));
 sg13g2_mux2_1 _10405_ (.A0(net3000),
    .A1(\cpu.regs[13][16] ),
    .S(net3225),
    .X(_00711_));
 sg13g2_a21oi_1 _10406_ (.A1(net3695),
    .A2(_03476_),
    .Y(_04699_),
    .B1(net3032));
 sg13g2_nor2_1 _10407_ (.A(_04041_),
    .B(net3376),
    .Y(_04700_));
 sg13g2_nor2_1 _10408_ (.A(net3310),
    .B(_04647_),
    .Y(_04701_));
 sg13g2_nand2b_1 _10409_ (.Y(_04702_),
    .B(_03856_),
    .A_N(_03854_));
 sg13g2_or2_1 _10410_ (.X(_04703_),
    .B(_04702_),
    .A(net3453));
 sg13g2_nand2_1 _10411_ (.Y(_04704_),
    .A(net3371),
    .B(_04702_));
 sg13g2_a22oi_1 _10412_ (.Y(_04705_),
    .B1(net3408),
    .B2(_04704_),
    .A2(_03857_),
    .A1(_03854_));
 sg13g2_o21ai_1 _10413_ (.B1(_04703_),
    .Y(_04706_),
    .A1(net3340),
    .A2(_04651_));
 sg13g2_nor4_2 _10414_ (.A(_04700_),
    .B(_04701_),
    .C(_04705_),
    .Y(_04707_),
    .D(_04706_));
 sg13g2_a22oi_1 _10415_ (.Y(_04708_),
    .B1(net3314),
    .B2(\cpu.PCreg0[17] ),
    .A2(net3381),
    .A1(\cpu.PC[17] ));
 sg13g2_o21ai_1 _10416_ (.B1(_04708_),
    .Y(_04709_),
    .A1(net3357),
    .A2(_04707_));
 sg13g2_nor2_2 _10417_ (.A(_04699_),
    .B(_04709_),
    .Y(_04710_));
 sg13g2_nand2_1 _10418_ (.Y(_04711_),
    .A(\cpu.regs[13][17] ),
    .B(net3223));
 sg13g2_o21ai_1 _10419_ (.B1(_04711_),
    .Y(_00712_),
    .A1(net3223),
    .A2(net2998));
 sg13g2_a21o_1 _10420_ (.A2(_03493_),
    .A1(net3697),
    .B1(net3031),
    .X(_04712_));
 sg13g2_nor2_1 _10421_ (.A(_03999_),
    .B(net3377),
    .Y(_04713_));
 sg13g2_nand2_1 _10422_ (.Y(_04714_),
    .A(_03847_),
    .B(_03849_));
 sg13g2_a21o_1 _10423_ (.A2(_04714_),
    .A1(net3371),
    .B1(net3410),
    .X(_04715_));
 sg13g2_o21ai_1 _10424_ (.B1(_04715_),
    .Y(_04716_),
    .A1(_03847_),
    .A2(_03849_));
 sg13g2_o21ai_1 _10425_ (.B1(_04716_),
    .Y(_04717_),
    .A1(net3453),
    .A2(_04714_));
 sg13g2_a21oi_1 _10426_ (.A1(net3312),
    .A2(_04626_),
    .Y(_04718_),
    .B1(_04717_));
 sg13g2_o21ai_1 _10427_ (.B1(_04718_),
    .Y(_04719_),
    .A1(net3340),
    .A2(_04630_));
 sg13g2_o21ai_1 _10428_ (.B1(net3355),
    .Y(_04720_),
    .A1(_04713_),
    .A2(_04719_));
 sg13g2_a22oi_1 _10429_ (.Y(_04721_),
    .B1(net3316),
    .B2(\cpu.PCreg0[18] ),
    .A2(net3379),
    .A1(\cpu.PC[18] ));
 sg13g2_nand3_1 _10430_ (.B(_04720_),
    .C(_04721_),
    .A(_04712_),
    .Y(_04722_));
 sg13g2_mux2_1 _10431_ (.A0(net2996),
    .A1(\cpu.regs[13][18] ),
    .S(net3224),
    .X(_00713_));
 sg13g2_a21oi_1 _10432_ (.A1(net3697),
    .A2(_03502_),
    .Y(_04723_),
    .B1(net3031));
 sg13g2_nor2_1 _10433_ (.A(net3343),
    .B(_04609_),
    .Y(_04724_));
 sg13g2_nand2b_1 _10434_ (.Y(_04725_),
    .B(_03839_),
    .A_N(_03837_));
 sg13g2_nand2_1 _10435_ (.Y(_04726_),
    .A(net3373),
    .B(_04725_));
 sg13g2_a22oi_1 _10436_ (.Y(_04727_),
    .B1(net3408),
    .B2(_04726_),
    .A2(_03840_),
    .A1(_03837_));
 sg13g2_nor2_1 _10437_ (.A(net3452),
    .B(_04725_),
    .Y(_04728_));
 sg13g2_nor3_1 _10438_ (.A(_04724_),
    .B(_04727_),
    .C(_04728_),
    .Y(_04729_));
 sg13g2_o21ai_1 _10439_ (.B1(_04729_),
    .Y(_04730_),
    .A1(_04008_),
    .A2(net3376));
 sg13g2_a21oi_1 _10440_ (.A1(net3312),
    .A2(_04605_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_a22oi_1 _10441_ (.Y(_04732_),
    .B1(net3318),
    .B2(\cpu.PCreg0[19] ),
    .A2(net3380),
    .A1(\cpu.PC[19] ));
 sg13g2_o21ai_1 _10442_ (.B1(_04732_),
    .Y(_04733_),
    .A1(net3357),
    .A2(_04731_));
 sg13g2_nor2_2 _10443_ (.A(_04723_),
    .B(_04733_),
    .Y(_04734_));
 sg13g2_nand2_1 _10444_ (.Y(_04735_),
    .A(\cpu.regs[13][19] ),
    .B(net3223));
 sg13g2_o21ai_1 _10445_ (.B1(_04735_),
    .Y(_00714_),
    .A1(net3223),
    .A2(net2994));
 sg13g2_a21oi_2 _10446_ (.B1(net3032),
    .Y(_04736_),
    .A2(_03516_),
    .A1(net3698));
 sg13g2_nor2_1 _10447_ (.A(_04004_),
    .B(net3376),
    .Y(_04737_));
 sg13g2_and3_1 _10448_ (.X(_04738_),
    .A(net3359),
    .B(_03871_),
    .C(_03872_));
 sg13g2_nor2b_1 _10449_ (.A(_03871_),
    .B_N(_03873_),
    .Y(_04739_));
 sg13g2_nand2b_1 _10450_ (.Y(_04740_),
    .B(net3371),
    .A_N(_04739_));
 sg13g2_a21oi_1 _10451_ (.A1(net3409),
    .A2(_04740_),
    .Y(_04741_),
    .B1(_04738_));
 sg13g2_a221oi_1 _10452_ (.B2(_04253_),
    .C1(_04741_),
    .B1(_04739_),
    .A1(net3312),
    .Y(_04742_),
    .A2(_04580_));
 sg13g2_o21ai_1 _10453_ (.B1(_04742_),
    .Y(_04743_),
    .A1(net3343),
    .A2(_04587_));
 sg13g2_o21ai_1 _10454_ (.B1(net3356),
    .Y(_04744_),
    .A1(_04737_),
    .A2(_04743_));
 sg13g2_a22oi_1 _10455_ (.Y(_04745_),
    .B1(net3315),
    .B2(\cpu.PCreg0[20] ),
    .A2(net3379),
    .A1(\cpu.PC[20] ));
 sg13g2_nand3b_1 _10456_ (.B(_04744_),
    .C(_04745_),
    .Y(_04746_),
    .A_N(_04736_));
 sg13g2_mux2_1 _10457_ (.A0(net2992),
    .A1(\cpu.regs[13][20] ),
    .S(net3220),
    .X(_00715_));
 sg13g2_a21o_1 _10458_ (.A2(_03529_),
    .A1(net3696),
    .B1(net3032),
    .X(_04747_));
 sg13g2_nand2_1 _10459_ (.Y(_04748_),
    .A(_03864_),
    .B(_03866_));
 sg13g2_a21o_1 _10460_ (.A2(_04748_),
    .A1(net3371),
    .B1(net3410),
    .X(_04749_));
 sg13g2_o21ai_1 _10461_ (.B1(_04749_),
    .Y(_04750_),
    .A1(_03864_),
    .A2(_03866_));
 sg13g2_o21ai_1 _10462_ (.B1(_04750_),
    .Y(_04751_),
    .A1(net3453),
    .A2(_04748_));
 sg13g2_a21o_1 _10463_ (.A2(_04552_),
    .A1(net3312),
    .B1(_04751_),
    .X(_04752_));
 sg13g2_nand2_1 _10464_ (.Y(_04753_),
    .A(net3348),
    .B(_04561_));
 sg13g2_o21ai_1 _10465_ (.B1(_04753_),
    .Y(_04754_),
    .A1(_04009_),
    .A2(net3376));
 sg13g2_o21ai_1 _10466_ (.B1(net3355),
    .Y(_04755_),
    .A1(_04752_),
    .A2(_04754_));
 sg13g2_a22oi_1 _10467_ (.Y(_04756_),
    .B1(net3316),
    .B2(\cpu.PCreg0[21] ),
    .A2(net3379),
    .A1(\cpu.PC[21] ));
 sg13g2_nand3_1 _10468_ (.B(_04755_),
    .C(_04756_),
    .A(_04747_),
    .Y(_04757_));
 sg13g2_mux2_1 _10469_ (.A0(net2990),
    .A1(\cpu.regs[13][21] ),
    .S(net3224),
    .X(_00716_));
 sg13g2_nor2_2 _10470_ (.A(net3624),
    .B(\cdi[22] ),
    .Y(_04758_));
 sg13g2_and3_1 _10471_ (.X(_04759_),
    .A(net3359),
    .B(_03888_),
    .C(_03889_));
 sg13g2_nor2b_1 _10472_ (.A(_03888_),
    .B_N(_03890_),
    .Y(_04760_));
 sg13g2_nand2b_1 _10473_ (.Y(_04761_),
    .B(net3372),
    .A_N(_04760_));
 sg13g2_a21oi_1 _10474_ (.A1(net3408),
    .A2(_04761_),
    .Y(_04762_),
    .B1(_04759_));
 sg13g2_a221oi_1 _10475_ (.B2(_04253_),
    .C1(_04762_),
    .B1(_04760_),
    .A1(net3312),
    .Y(_04763_),
    .A2(_04523_));
 sg13g2_o21ai_1 _10476_ (.B1(_04763_),
    .Y(_04764_),
    .A1(net3343),
    .A2(_04532_));
 sg13g2_a21oi_1 _10477_ (.A1(_04012_),
    .A2(net3337),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nor2_1 _10478_ (.A(net3357),
    .B(_04765_),
    .Y(_04766_));
 sg13g2_a221oi_1 _10479_ (.B2(\cpu.PCreg0[22] ),
    .C1(_04766_),
    .B1(net3316),
    .A1(\cpu.PC[22] ),
    .Y(_04767_),
    .A2(net3379));
 sg13g2_o21ai_1 _10480_ (.B1(_04767_),
    .Y(_04768_),
    .A1(net3031),
    .A2(_04758_));
 sg13g2_mux2_1 _10481_ (.A0(net3017),
    .A1(\cpu.regs[13][22] ),
    .S(net3221),
    .X(_00717_));
 sg13g2_nor2_2 _10482_ (.A(net3624),
    .B(\cdi[23] ),
    .Y(_04769_));
 sg13g2_nor2_1 _10483_ (.A(_03983_),
    .B(net3376),
    .Y(_04770_));
 sg13g2_nand2_1 _10484_ (.Y(_04771_),
    .A(_03896_),
    .B(_03898_));
 sg13g2_a21o_1 _10485_ (.A2(_04771_),
    .A1(net3371),
    .B1(net3410),
    .X(_04772_));
 sg13g2_o21ai_1 _10486_ (.B1(_04772_),
    .Y(_04773_),
    .A1(_03896_),
    .A2(_03898_));
 sg13g2_o21ai_1 _10487_ (.B1(_04773_),
    .Y(_04774_),
    .A1(net3452),
    .A2(_04771_));
 sg13g2_a21oi_1 _10488_ (.A1(net3312),
    .A2(_04500_),
    .Y(_04775_),
    .B1(_04774_));
 sg13g2_o21ai_1 _10489_ (.B1(_04775_),
    .Y(_04776_),
    .A1(net3343),
    .A2(_04510_));
 sg13g2_o21ai_1 _10490_ (.B1(net3355),
    .Y(_04777_),
    .A1(_04770_),
    .A2(_04776_));
 sg13g2_a22oi_1 _10491_ (.Y(_04778_),
    .B1(net3316),
    .B2(\cpu.PCreg0[23] ),
    .A2(net3380),
    .A1(\cpu.PC[23] ));
 sg13g2_and2_1 _10492_ (.A(_04777_),
    .B(_04778_),
    .X(_04779_));
 sg13g2_o21ai_1 _10493_ (.B1(_04779_),
    .Y(_04780_),
    .A1(net3031),
    .A2(_04769_));
 sg13g2_mux2_1 _10494_ (.A0(net3016),
    .A1(\cpu.regs[13][23] ),
    .S(net3221),
    .X(_00718_));
 sg13g2_a21o_1 _10495_ (.A2(_03573_),
    .A1(net3696),
    .B1(net3032),
    .X(_04781_));
 sg13g2_or2_1 _10496_ (.X(_04782_),
    .B(_03937_),
    .A(_03936_));
 sg13g2_a21oi_1 _10497_ (.A1(net3375),
    .A2(_04782_),
    .Y(_04783_),
    .B1(net3412));
 sg13g2_a21o_1 _10498_ (.A2(_03937_),
    .A1(_03936_),
    .B1(_04783_),
    .X(_04784_));
 sg13g2_o21ai_1 _10499_ (.B1(_04784_),
    .Y(_04785_),
    .A1(net3455),
    .A2(_04782_));
 sg13g2_a221oi_1 _10500_ (.B2(net3313),
    .C1(_04785_),
    .B1(_04478_),
    .A1(net3352),
    .Y(_04786_),
    .A2(_04472_));
 sg13g2_o21ai_1 _10501_ (.B1(_04786_),
    .Y(_04787_),
    .A1(_04039_),
    .A2(net3376));
 sg13g2_nand2_1 _10502_ (.Y(_04788_),
    .A(net3356),
    .B(_04787_));
 sg13g2_a22oi_1 _10503_ (.Y(_04789_),
    .B1(net3316),
    .B2(\cpu.PCreg0[24] ),
    .A2(net3379),
    .A1(\cpu.PC[24] ));
 sg13g2_nand3_1 _10504_ (.B(_04788_),
    .C(_04789_),
    .A(_04781_),
    .Y(_04790_));
 sg13g2_mux2_1 _10505_ (.A0(net2987),
    .A1(\cpu.regs[13][24] ),
    .S(net3221),
    .X(_00719_));
 sg13g2_a21o_1 _10506_ (.A2(_03581_),
    .A1(net3696),
    .B1(net3032),
    .X(_04791_));
 sg13g2_nor2_1 _10507_ (.A(_04045_),
    .B(net3376),
    .Y(_04792_));
 sg13g2_or2_1 _10508_ (.X(_04793_),
    .B(_03931_),
    .A(_03930_));
 sg13g2_a21oi_1 _10509_ (.A1(net3375),
    .A2(_04793_),
    .Y(_04794_),
    .B1(net3411));
 sg13g2_a21o_1 _10510_ (.A2(_03931_),
    .A1(_03930_),
    .B1(_04794_),
    .X(_04795_));
 sg13g2_o21ai_1 _10511_ (.B1(_04795_),
    .Y(_04796_),
    .A1(net3455),
    .A2(_04793_));
 sg13g2_a21oi_1 _10512_ (.A1(_04264_),
    .A2(_04431_),
    .Y(_04797_),
    .B1(_04796_));
 sg13g2_o21ai_1 _10513_ (.B1(_04797_),
    .Y(_04798_),
    .A1(net3344),
    .A2(_04440_));
 sg13g2_o21ai_1 _10514_ (.B1(net3355),
    .Y(_04799_),
    .A1(_04792_),
    .A2(_04798_));
 sg13g2_a22oi_1 _10515_ (.Y(_04800_),
    .B1(net3316),
    .B2(\cpu.PCreg0[25] ),
    .A2(net3380),
    .A1(\cpu.PC[25] ));
 sg13g2_nand3_1 _10516_ (.B(_04799_),
    .C(_04800_),
    .A(_04791_),
    .Y(_04801_));
 sg13g2_mux2_1 _10517_ (.A0(net2986),
    .A1(\cpu.regs[13][25] ),
    .S(net3224),
    .X(_00720_));
 sg13g2_nor2_2 _10518_ (.A(net3624),
    .B(\cdi[26] ),
    .Y(_04802_));
 sg13g2_nor2_1 _10519_ (.A(_03923_),
    .B(_03926_),
    .Y(_04803_));
 sg13g2_o21ai_1 _10520_ (.B1(net3371),
    .Y(_04804_),
    .A1(_03923_),
    .A2(_03926_));
 sg13g2_a22oi_1 _10521_ (.Y(_04805_),
    .B1(net3408),
    .B2(_04804_),
    .A2(_03926_),
    .A1(_03923_));
 sg13g2_a221oi_1 _10522_ (.B2(_04253_),
    .C1(_04805_),
    .B1(_04803_),
    .A1(net3312),
    .Y(_04806_),
    .A2(_04397_));
 sg13g2_a22oi_1 _10523_ (.Y(_04807_),
    .B1(_04411_),
    .B2(net3348),
    .A2(net3337),
    .A1(_03995_));
 sg13g2_a21oi_2 _10524_ (.B1(net3357),
    .Y(_04808_),
    .A2(_04807_),
    .A1(_04806_));
 sg13g2_a221oi_1 _10525_ (.B2(\cpu.PCreg0[26] ),
    .C1(_04808_),
    .B1(net3316),
    .A1(\cpu.PC[26] ),
    .Y(_04809_),
    .A2(net3380));
 sg13g2_o21ai_1 _10526_ (.B1(_04809_),
    .Y(_04810_),
    .A1(net3031),
    .A2(_04802_));
 sg13g2_mux2_1 _10527_ (.A0(net3014),
    .A1(\cpu.regs[13][26] ),
    .S(net3221),
    .X(_00721_));
 sg13g2_nor2_2 _10528_ (.A(net3625),
    .B(\cdi[27] ),
    .Y(_04811_));
 sg13g2_nor2_1 _10529_ (.A(_04011_),
    .B(net3376),
    .Y(_04812_));
 sg13g2_nor2_2 _10530_ (.A(net3311),
    .B(_04379_),
    .Y(_04813_));
 sg13g2_nor2_2 _10531_ (.A(net3347),
    .B(_04370_),
    .Y(_04814_));
 sg13g2_nand2_1 _10532_ (.Y(_04815_),
    .A(_03916_),
    .B(_03919_));
 sg13g2_a21o_1 _10533_ (.A2(_04815_),
    .A1(net3371),
    .B1(net3410),
    .X(_04816_));
 sg13g2_o21ai_1 _10534_ (.B1(_04816_),
    .Y(_04817_),
    .A1(_03916_),
    .A2(_03919_));
 sg13g2_o21ai_1 _10535_ (.B1(_04817_),
    .Y(_04818_),
    .A1(net3452),
    .A2(_04815_));
 sg13g2_nor4_1 _10536_ (.A(_04812_),
    .B(_04813_),
    .C(_04814_),
    .D(_04818_),
    .Y(_04819_));
 sg13g2_nor2_1 _10537_ (.A(net3357),
    .B(_04819_),
    .Y(_04820_));
 sg13g2_a221oi_1 _10538_ (.B2(\cpu.PCreg0[27] ),
    .C1(_04820_),
    .B1(net3315),
    .A1(\cpu.PC[27] ),
    .Y(_04821_),
    .A2(net3379));
 sg13g2_o21ai_1 _10539_ (.B1(_04821_),
    .Y(_04822_),
    .A1(net3031),
    .A2(_04811_));
 sg13g2_mux2_1 _10540_ (.A0(net3012),
    .A1(\cpu.regs[13][27] ),
    .S(net3221),
    .X(_00722_));
 sg13g2_a21o_1 _10541_ (.A2(_03595_),
    .A1(net3695),
    .B1(net3032),
    .X(_04823_));
 sg13g2_nor2_1 _10542_ (.A(_04015_),
    .B(net3377),
    .Y(_04824_));
 sg13g2_nand2_1 _10543_ (.Y(_04825_),
    .A(_03957_),
    .B(_03959_));
 sg13g2_a21o_1 _10544_ (.A2(_04825_),
    .A1(net3373),
    .B1(net3410),
    .X(_04826_));
 sg13g2_o21ai_1 _10545_ (.B1(_04826_),
    .Y(_04827_),
    .A1(_03957_),
    .A2(_03959_));
 sg13g2_o21ai_1 _10546_ (.B1(_04827_),
    .Y(_04828_),
    .A1(net3452),
    .A2(_04825_));
 sg13g2_a21oi_1 _10547_ (.A1(net3313),
    .A2(_04345_),
    .Y(_04829_),
    .B1(_04828_));
 sg13g2_o21ai_1 _10548_ (.B1(_04829_),
    .Y(_04830_),
    .A1(net3345),
    .A2(_04337_));
 sg13g2_o21ai_1 _10549_ (.B1(net3355),
    .Y(_04831_),
    .A1(_04824_),
    .A2(_04830_));
 sg13g2_a22oi_1 _10550_ (.Y(_04832_),
    .B1(net3315),
    .B2(\cpu.PCreg0[28] ),
    .A2(net3379),
    .A1(\cpu.PC[28] ));
 sg13g2_nand3_1 _10551_ (.B(_04831_),
    .C(_04832_),
    .A(_04823_),
    .Y(_04833_));
 sg13g2_mux2_1 _10552_ (.A0(net2983),
    .A1(\cpu.regs[13][28] ),
    .S(net3221),
    .X(_00723_));
 sg13g2_a21o_1 _10553_ (.A2(_03599_),
    .A1(net3698),
    .B1(net3032),
    .X(_04834_));
 sg13g2_nand2_1 _10554_ (.Y(_04835_),
    .A(_03950_),
    .B(_03952_));
 sg13g2_a21o_1 _10555_ (.A2(_04835_),
    .A1(net3374),
    .B1(net3411),
    .X(_04836_));
 sg13g2_o21ai_1 _10556_ (.B1(_04836_),
    .Y(_04837_),
    .A1(_03950_),
    .A2(_03952_));
 sg13g2_o21ai_1 _10557_ (.B1(_04837_),
    .Y(_04838_),
    .A1(net3454),
    .A2(_04835_));
 sg13g2_a221oi_1 _10558_ (.B2(net3353),
    .C1(_04838_),
    .B1(_04317_),
    .A1(net3313),
    .Y(_04839_),
    .A2(_04308_));
 sg13g2_o21ai_1 _10559_ (.B1(_04839_),
    .Y(_04840_),
    .A1(_04048_),
    .A2(net3377));
 sg13g2_nand2_1 _10560_ (.Y(_04841_),
    .A(net3355),
    .B(_04840_));
 sg13g2_a22oi_1 _10561_ (.Y(_04842_),
    .B1(net3314),
    .B2(\cpu.PCreg0[29] ),
    .A2(net3381),
    .A1(\cpu.PC[29] ));
 sg13g2_nand3_1 _10562_ (.B(_04841_),
    .C(_04842_),
    .A(_04834_),
    .Y(_04843_));
 sg13g2_mux2_1 _10563_ (.A0(net2982),
    .A1(\cpu.regs[13][29] ),
    .S(net3221),
    .X(_00724_));
 sg13g2_nor2_1 _10564_ (.A(net3625),
    .B(\cdi[30] ),
    .Y(_04844_));
 sg13g2_nand2_1 _10565_ (.Y(_04845_),
    .A(_03666_),
    .B(_03670_));
 sg13g2_a21o_1 _10566_ (.A2(_04845_),
    .A1(net3373),
    .B1(net3410),
    .X(_04846_));
 sg13g2_o21ai_1 _10567_ (.B1(_04846_),
    .Y(_04847_),
    .A1(_03666_),
    .A2(_03670_));
 sg13g2_o21ai_1 _10568_ (.B1(_04847_),
    .Y(_04848_),
    .A1(net3452),
    .A2(_04845_));
 sg13g2_a21oi_1 _10569_ (.A1(net3312),
    .A2(_04282_),
    .Y(_04849_),
    .B1(_04848_));
 sg13g2_nor2_2 _10570_ (.A(net3347),
    .B(_04274_),
    .Y(_04850_));
 sg13g2_a21oi_1 _10571_ (.A1(_04014_),
    .A2(net3337),
    .Y(_04851_),
    .B1(_04850_));
 sg13g2_a21oi_1 _10572_ (.A1(_04849_),
    .A2(_04851_),
    .Y(_04852_),
    .B1(net3357));
 sg13g2_a221oi_1 _10573_ (.B2(\cpu.PCreg0[30] ),
    .C1(_04852_),
    .B1(net3314),
    .A1(\cpu.PC[30] ),
    .Y(_04853_),
    .A2(net3381));
 sg13g2_o21ai_1 _10574_ (.B1(_04853_),
    .Y(_04854_),
    .A1(net3031),
    .A2(_04844_));
 sg13g2_mux2_1 _10575_ (.A0(net3009),
    .A1(\cpu.regs[13][30] ),
    .S(net3220),
    .X(_00725_));
 sg13g2_nor2_1 _10576_ (.A(net3625),
    .B(\cdi[31] ),
    .Y(_04855_));
 sg13g2_nor2_1 _10577_ (.A(net3347),
    .B(_04231_),
    .Y(_04856_));
 sg13g2_nor2_1 _10578_ (.A(_04247_),
    .B(net3311),
    .Y(_04857_));
 sg13g2_nand2b_1 _10579_ (.Y(_04858_),
    .B(net3374),
    .A_N(_03972_));
 sg13g2_nand3_1 _10580_ (.B(_03661_),
    .C(_04253_),
    .A(_03657_),
    .Y(_04859_));
 sg13g2_o21ai_1 _10581_ (.B1(net3411),
    .Y(_04860_),
    .A1(_03657_),
    .A2(_03661_));
 sg13g2_nand3_1 _10582_ (.B(_04859_),
    .C(_04860_),
    .A(_04858_),
    .Y(_04861_));
 sg13g2_nor3_2 _10583_ (.A(_04856_),
    .B(_04857_),
    .C(_04861_),
    .Y(_04862_));
 sg13g2_o21ai_1 _10584_ (.B1(_04862_),
    .Y(_04863_),
    .A1(_04013_),
    .A2(net3377));
 sg13g2_and2_1 _10585_ (.A(\cpu.PC[31] ),
    .B(net3379),
    .X(_04864_));
 sg13g2_a221oi_1 _10586_ (.B2(net3355),
    .C1(_04864_),
    .B1(_04863_),
    .A1(\cpu.PCreg0[31] ),
    .Y(_04865_),
    .A2(net3315));
 sg13g2_o21ai_1 _10587_ (.B1(_04865_),
    .Y(_04866_),
    .A1(net3031),
    .A2(_04855_));
 sg13g2_mux2_1 _10588_ (.A0(net3008),
    .A1(\cpu.regs[13][31] ),
    .S(net3221),
    .X(_00726_));
 sg13g2_nand2_1 _10589_ (.Y(_04867_),
    .A(net3098),
    .B(_03425_));
 sg13g2_nand4_1 _10590_ (.B(net3450),
    .C(net3099),
    .A(net3698),
    .Y(_04868_),
    .D(_03425_));
 sg13g2_nor3_2 _10591_ (.A(net3125),
    .B(_03442_),
    .C(_04868_),
    .Y(_04869_));
 sg13g2_mux2_1 _10592_ (.A0(\irqvect[1][0] ),
    .A1(net3326),
    .S(net3083),
    .X(_00727_));
 sg13g2_mux2_1 _10593_ (.A0(\irqvect[1][1] ),
    .A1(net3327),
    .S(net3084),
    .X(_00728_));
 sg13g2_nor2_1 _10594_ (.A(\irqvect[1][2] ),
    .B(net3083),
    .Y(_04870_));
 sg13g2_a21oi_1 _10595_ (.A1(_02928_),
    .A2(net3083),
    .Y(_00729_),
    .B1(_04870_));
 sg13g2_mux2_1 _10596_ (.A0(\irqvect[1][3] ),
    .A1(net3328),
    .S(net3084),
    .X(_00730_));
 sg13g2_mux2_1 _10597_ (.A0(\irqvect[1][4] ),
    .A1(net3329),
    .S(net3084),
    .X(_00731_));
 sg13g2_mux2_1 _10598_ (.A0(\irqvect[1][5] ),
    .A1(net3330),
    .S(net3084),
    .X(_00732_));
 sg13g2_nor2_1 _10599_ (.A(\irqvect[1][6] ),
    .B(net3084),
    .Y(_04871_));
 sg13g2_a21oi_1 _10600_ (.A1(_03267_),
    .A2(net3084),
    .Y(_00733_),
    .B1(_04871_));
 sg13g2_nor2_1 _10601_ (.A(\irqvect[1][7] ),
    .B(net3084),
    .Y(_04872_));
 sg13g2_a21oi_1 _10602_ (.A1(_03193_),
    .A2(net3084),
    .Y(_00734_),
    .B1(_04872_));
 sg13g2_nor2_1 _10603_ (.A(\irqvect[1][8] ),
    .B(net3085),
    .Y(_04873_));
 sg13g2_a21oi_1 _10604_ (.A1(_03120_),
    .A2(net3085),
    .Y(_00735_),
    .B1(_04873_));
 sg13g2_nor2_1 _10605_ (.A(\irqvect[1][9] ),
    .B(net3080),
    .Y(_04874_));
 sg13g2_a21oi_1 _10606_ (.A1(_03033_),
    .A2(net3080),
    .Y(_00736_),
    .B1(_04874_));
 sg13g2_nor2_1 _10607_ (.A(\irqvect[1][10] ),
    .B(net3085),
    .Y(_04875_));
 sg13g2_a21oi_1 _10608_ (.A1(_02947_),
    .A2(net3083),
    .Y(_00737_),
    .B1(_04875_));
 sg13g2_nor2_1 _10609_ (.A(\irqvect[1][11] ),
    .B(net3082),
    .Y(_04876_));
 sg13g2_a21oi_1 _10610_ (.A1(_02861_),
    .A2(net3082),
    .Y(_00738_),
    .B1(_04876_));
 sg13g2_nor2_1 _10611_ (.A(\irqvect[1][12] ),
    .B(net3081),
    .Y(_04877_));
 sg13g2_a21oi_1 _10612_ (.A1(_02778_),
    .A2(net3081),
    .Y(_00739_),
    .B1(_04877_));
 sg13g2_nor2_1 _10613_ (.A(\irqvect[1][13] ),
    .B(_04869_),
    .Y(_04878_));
 sg13g2_a21oi_1 _10614_ (.A1(_02682_),
    .A2(net3085),
    .Y(_00740_),
    .B1(_04878_));
 sg13g2_nor2_1 _10615_ (.A(\irqvect[1][14] ),
    .B(net3083),
    .Y(_04879_));
 sg13g2_a21oi_1 _10616_ (.A1(_03288_),
    .A2(net3083),
    .Y(_00741_),
    .B1(_04879_));
 sg13g2_nor2_1 _10617_ (.A(\irqvect[1][15] ),
    .B(net3083),
    .Y(_04880_));
 sg13g2_a21oi_1 _10618_ (.A1(_03216_),
    .A2(net3083),
    .Y(_00742_),
    .B1(_04880_));
 sg13g2_nor2_1 _10619_ (.A(\irqvect[1][16] ),
    .B(net3078),
    .Y(_04881_));
 sg13g2_a21oi_1 _10620_ (.A1(_03142_),
    .A2(net3078),
    .Y(_00743_),
    .B1(_04881_));
 sg13g2_nor2_1 _10621_ (.A(\irqvect[1][17] ),
    .B(net3079),
    .Y(_04882_));
 sg13g2_a21oi_1 _10622_ (.A1(_03054_),
    .A2(net3079),
    .Y(_00744_),
    .B1(_04882_));
 sg13g2_nor2_1 _10623_ (.A(\irqvect[1][18] ),
    .B(net3079),
    .Y(_04883_));
 sg13g2_a21oi_1 _10624_ (.A1(_02967_),
    .A2(net3079),
    .Y(_00745_),
    .B1(_04883_));
 sg13g2_nor2_1 _10625_ (.A(\irqvect[1][19] ),
    .B(net3078),
    .Y(_04884_));
 sg13g2_a21oi_1 _10626_ (.A1(_02881_),
    .A2(net3078),
    .Y(_00746_),
    .B1(_04884_));
 sg13g2_nor2_1 _10627_ (.A(\irqvect[1][20] ),
    .B(net3079),
    .Y(_04885_));
 sg13g2_a21oi_1 _10628_ (.A1(_02798_),
    .A2(net3079),
    .Y(_00747_),
    .B1(_04885_));
 sg13g2_nor2_1 _10629_ (.A(\irqvect[1][21] ),
    .B(net3081),
    .Y(_04886_));
 sg13g2_a21oi_1 _10630_ (.A1(_02703_),
    .A2(net3081),
    .Y(_00748_),
    .B1(_04886_));
 sg13g2_nor2_1 _10631_ (.A(\irqvect[1][22] ),
    .B(net3080),
    .Y(_04887_));
 sg13g2_a21oi_1 _10632_ (.A1(_03269_),
    .A2(net3080),
    .Y(_00749_),
    .B1(_04887_));
 sg13g2_nor2_1 _10633_ (.A(\irqvect[1][23] ),
    .B(net3080),
    .Y(_04888_));
 sg13g2_a21oi_1 _10634_ (.A1(_03195_),
    .A2(net3080),
    .Y(_00750_),
    .B1(_04888_));
 sg13g2_nor2_1 _10635_ (.A(\irqvect[1][24] ),
    .B(net3080),
    .Y(_04889_));
 sg13g2_a21oi_1 _10636_ (.A1(_03122_),
    .A2(net3080),
    .Y(_00751_),
    .B1(_04889_));
 sg13g2_nor2_1 _10637_ (.A(\irqvect[1][25] ),
    .B(net3085),
    .Y(_04890_));
 sg13g2_a21oi_1 _10638_ (.A1(_03035_),
    .A2(net3085),
    .Y(_00752_),
    .B1(_04890_));
 sg13g2_nor2_1 _10639_ (.A(\irqvect[1][26] ),
    .B(net3079),
    .Y(_04891_));
 sg13g2_a21oi_1 _10640_ (.A1(_02949_),
    .A2(net3079),
    .Y(_00753_),
    .B1(_04891_));
 sg13g2_nor2_1 _10641_ (.A(\irqvect[1][27] ),
    .B(net3081),
    .Y(_04892_));
 sg13g2_a21oi_1 _10642_ (.A1(_02863_),
    .A2(net3081),
    .Y(_00754_),
    .B1(_04892_));
 sg13g2_nor2_1 _10643_ (.A(\irqvect[1][28] ),
    .B(net3078),
    .Y(_04893_));
 sg13g2_a21oi_1 _10644_ (.A1(_02780_),
    .A2(net3078),
    .Y(_00755_),
    .B1(_04893_));
 sg13g2_nor2_1 _10645_ (.A(\irqvect[1][29] ),
    .B(net3078),
    .Y(_04894_));
 sg13g2_a21oi_1 _10646_ (.A1(_02684_),
    .A2(net3078),
    .Y(_00756_),
    .B1(_04894_));
 sg13g2_nand2_1 _10647_ (.Y(_04895_),
    .A(\cpu.Bimm[2] ),
    .B(net3701));
 sg13g2_nand2_1 _10648_ (.Y(_04896_),
    .A(_04123_),
    .B(_04895_));
 sg13g2_nor2_1 _10649_ (.A(_04122_),
    .B(_04896_),
    .Y(_04897_));
 sg13g2_nand2_2 _10650_ (.Y(_04898_),
    .A(_04113_),
    .B(_04897_));
 sg13g2_mux2_1 _10651_ (.A0(net3046),
    .A1(\cpu.regs[1][0] ),
    .S(net3219),
    .X(_00757_));
 sg13g2_mux2_1 _10652_ (.A0(net3041),
    .A1(\cpu.regs[1][1] ),
    .S(net3219),
    .X(_00758_));
 sg13g2_mux2_1 _10653_ (.A0(net3040),
    .A1(\cpu.regs[1][2] ),
    .S(net3219),
    .X(_00759_));
 sg13g2_mux2_1 _10654_ (.A0(net3005),
    .A1(\cpu.regs[1][3] ),
    .S(net3218),
    .X(_00760_));
 sg13g2_mux2_1 _10655_ (.A0(net3003),
    .A1(\cpu.regs[1][4] ),
    .S(net3219),
    .X(_00761_));
 sg13g2_mux2_1 _10656_ (.A0(net3029),
    .A1(\cpu.regs[1][5] ),
    .S(net3218),
    .X(_00762_));
 sg13g2_mux2_1 _10657_ (.A0(net3037),
    .A1(\cpu.regs[1][6] ),
    .S(net3219),
    .X(_00763_));
 sg13g2_mux2_1 _10658_ (.A0(net3044),
    .A1(\cpu.regs[1][7] ),
    .S(net3218),
    .X(_00764_));
 sg13g2_mux2_1 _10659_ (.A0(net3027),
    .A1(\cpu.regs[1][8] ),
    .S(net3218),
    .X(_00765_));
 sg13g2_mux2_1 _10660_ (.A0(net3026),
    .A1(\cpu.regs[1][9] ),
    .S(net3217),
    .X(_00766_));
 sg13g2_mux2_1 _10661_ (.A0(net3023),
    .A1(\cpu.regs[1][10] ),
    .S(net3218),
    .X(_00767_));
 sg13g2_mux2_1 _10662_ (.A0(net3021),
    .A1(\cpu.regs[1][11] ),
    .S(net3218),
    .X(_00768_));
 sg13g2_mux2_1 _10663_ (.A0(net3001),
    .A1(\cpu.regs[1][12] ),
    .S(net3216),
    .X(_00769_));
 sg13g2_mux2_1 _10664_ (.A0(net3019),
    .A1(\cpu.regs[1][13] ),
    .S(net3216),
    .X(_00770_));
 sg13g2_nand2_1 _10665_ (.Y(_04899_),
    .A(\cpu.regs[1][14] ),
    .B(net3217));
 sg13g2_o21ai_1 _10666_ (.B1(_04899_),
    .Y(_00771_),
    .A1(net3035),
    .A2(net3217));
 sg13g2_nand2_1 _10667_ (.Y(_04900_),
    .A(\cpu.regs[1][15] ),
    .B(net3217));
 sg13g2_o21ai_1 _10668_ (.B1(_04900_),
    .Y(_00772_),
    .A1(net3033),
    .A2(net3217));
 sg13g2_mux2_1 _10669_ (.A0(net2999),
    .A1(\cpu.regs[1][16] ),
    .S(net3219),
    .X(_00773_));
 sg13g2_nand2_1 _10670_ (.Y(_04901_),
    .A(\cpu.regs[1][17] ),
    .B(net3217));
 sg13g2_o21ai_1 _10671_ (.B1(_04901_),
    .Y(_00774_),
    .A1(net2997),
    .A2(net3217));
 sg13g2_mux2_1 _10672_ (.A0(net2995),
    .A1(\cpu.regs[1][18] ),
    .S(net3216),
    .X(_00775_));
 sg13g2_nand2_1 _10673_ (.Y(_04902_),
    .A(\cpu.regs[1][19] ),
    .B(net3218));
 sg13g2_o21ai_1 _10674_ (.B1(_04902_),
    .Y(_00776_),
    .A1(net2993),
    .A2(net3217));
 sg13g2_mux2_1 _10675_ (.A0(net2991),
    .A1(\cpu.regs[1][20] ),
    .S(net3216),
    .X(_00777_));
 sg13g2_mux2_1 _10676_ (.A0(net2990),
    .A1(\cpu.regs[1][21] ),
    .S(net3215),
    .X(_00778_));
 sg13g2_mux2_1 _10677_ (.A0(net3018),
    .A1(\cpu.regs[1][22] ),
    .S(net3215),
    .X(_00779_));
 sg13g2_mux2_1 _10678_ (.A0(net3015),
    .A1(\cpu.regs[1][23] ),
    .S(net3215),
    .X(_00780_));
 sg13g2_mux2_1 _10679_ (.A0(net2988),
    .A1(\cpu.regs[1][24] ),
    .S(net3215),
    .X(_00781_));
 sg13g2_mux2_1 _10680_ (.A0(net2985),
    .A1(\cpu.regs[1][25] ),
    .S(net3215),
    .X(_00782_));
 sg13g2_mux2_1 _10681_ (.A0(net3013),
    .A1(\cpu.regs[1][26] ),
    .S(net3216),
    .X(_00783_));
 sg13g2_mux2_1 _10682_ (.A0(net3011),
    .A1(\cpu.regs[1][27] ),
    .S(net3215),
    .X(_00784_));
 sg13g2_mux2_1 _10683_ (.A0(net2984),
    .A1(\cpu.regs[1][28] ),
    .S(net3215),
    .X(_00785_));
 sg13g2_mux2_1 _10684_ (.A0(net2981),
    .A1(\cpu.regs[1][29] ),
    .S(net3215),
    .X(_00786_));
 sg13g2_mux2_1 _10685_ (.A0(net3009),
    .A1(\cpu.regs[1][30] ),
    .S(net3216),
    .X(_00787_));
 sg13g2_mux2_1 _10686_ (.A0(net3007),
    .A1(\cpu.regs[1][31] ),
    .S(net3216),
    .X(_00788_));
 sg13g2_nand3_1 _10687_ (.B(\cpu.Bimm[11] ),
    .C(net3701),
    .A(\cpu.Bimm[1] ),
    .Y(_04903_));
 sg13g2_nor3_2 _10688_ (.A(\cpu.Bimm[2] ),
    .B(_04122_),
    .C(_04123_),
    .Y(_04904_));
 sg13g2_nor2b_1 _10689_ (.A(_04903_),
    .B_N(_04904_),
    .Y(_04905_));
 sg13g2_mux2_1 _10690_ (.A0(\cpu.regs[11][0] ),
    .A1(net3047),
    .S(net3213),
    .X(_00789_));
 sg13g2_mux2_1 _10691_ (.A0(\cpu.regs[11][1] ),
    .A1(net3041),
    .S(net3213),
    .X(_00790_));
 sg13g2_mux2_1 _10692_ (.A0(\cpu.regs[11][2] ),
    .A1(net3039),
    .S(net3213),
    .X(_00791_));
 sg13g2_mux2_1 _10693_ (.A0(\cpu.regs[11][3] ),
    .A1(net3006),
    .S(net3212),
    .X(_00792_));
 sg13g2_mux2_1 _10694_ (.A0(\cpu.regs[11][4] ),
    .A1(net3004),
    .S(net3213),
    .X(_00793_));
 sg13g2_mux2_1 _10695_ (.A0(\cpu.regs[11][5] ),
    .A1(net3030),
    .S(net3212),
    .X(_00794_));
 sg13g2_mux2_1 _10696_ (.A0(\cpu.regs[11][6] ),
    .A1(net3038),
    .S(net3213),
    .X(_00795_));
 sg13g2_mux2_1 _10697_ (.A0(\cpu.regs[11][7] ),
    .A1(net3045),
    .S(net3212),
    .X(_00796_));
 sg13g2_mux2_1 _10698_ (.A0(\cpu.regs[11][8] ),
    .A1(net3028),
    .S(net3212),
    .X(_00797_));
 sg13g2_mux2_1 _10699_ (.A0(\cpu.regs[11][9] ),
    .A1(net3025),
    .S(net3213),
    .X(_00798_));
 sg13g2_mux2_1 _10700_ (.A0(\cpu.regs[11][10] ),
    .A1(net3024),
    .S(net3211),
    .X(_00799_));
 sg13g2_mux2_1 _10701_ (.A0(\cpu.regs[11][11] ),
    .A1(net3022),
    .S(net3211),
    .X(_00800_));
 sg13g2_mux2_1 _10702_ (.A0(\cpu.regs[11][12] ),
    .A1(net3002),
    .S(net3210),
    .X(_00801_));
 sg13g2_mux2_1 _10703_ (.A0(\cpu.regs[11][13] ),
    .A1(net3020),
    .S(net3210),
    .X(_00802_));
 sg13g2_nor2_1 _10704_ (.A(\cpu.regs[11][14] ),
    .B(net3211),
    .Y(_04906_));
 sg13g2_a21oi_1 _10705_ (.A1(net3036),
    .A2(net3211),
    .Y(_00803_),
    .B1(_04906_));
 sg13g2_nor2_1 _10706_ (.A(\cpu.regs[11][15] ),
    .B(net3211),
    .Y(_04907_));
 sg13g2_a21oi_1 _10707_ (.A1(net3034),
    .A2(net3211),
    .Y(_00804_),
    .B1(_04907_));
 sg13g2_mux2_1 _10708_ (.A0(\cpu.regs[11][16] ),
    .A1(net3000),
    .S(net3213),
    .X(_00805_));
 sg13g2_nor2_1 _10709_ (.A(\cpu.regs[11][17] ),
    .B(net3211),
    .Y(_04908_));
 sg13g2_a21oi_1 _10710_ (.A1(net2998),
    .A2(net3211),
    .Y(_00806_),
    .B1(_04908_));
 sg13g2_mux2_1 _10711_ (.A0(\cpu.regs[11][18] ),
    .A1(net2996),
    .S(net3214),
    .X(_00807_));
 sg13g2_nor2_1 _10712_ (.A(\cpu.regs[11][19] ),
    .B(net3209),
    .Y(_04909_));
 sg13g2_a21oi_1 _10713_ (.A1(net2994),
    .A2(net3209),
    .Y(_00808_),
    .B1(_04909_));
 sg13g2_mux2_1 _10714_ (.A0(\cpu.regs[11][20] ),
    .A1(net2992),
    .S(net3210),
    .X(_00809_));
 sg13g2_mux2_1 _10715_ (.A0(\cpu.regs[11][21] ),
    .A1(net2990),
    .S(net3209),
    .X(_00810_));
 sg13g2_mux2_1 _10716_ (.A0(\cpu.regs[11][22] ),
    .A1(net3017),
    .S(net3209),
    .X(_00811_));
 sg13g2_mux2_1 _10717_ (.A0(\cpu.regs[11][23] ),
    .A1(net3016),
    .S(net3209),
    .X(_00812_));
 sg13g2_mux2_1 _10718_ (.A0(\cpu.regs[11][24] ),
    .A1(net2987),
    .S(net3209),
    .X(_00813_));
 sg13g2_mux2_1 _10719_ (.A0(\cpu.regs[11][25] ),
    .A1(net2986),
    .S(net3214),
    .X(_00814_));
 sg13g2_mux2_1 _10720_ (.A0(\cpu.regs[11][26] ),
    .A1(net3013),
    .S(net3210),
    .X(_00815_));
 sg13g2_mux2_1 _10721_ (.A0(\cpu.regs[11][27] ),
    .A1(net3012),
    .S(net3209),
    .X(_00816_));
 sg13g2_mux2_1 _10722_ (.A0(\cpu.regs[11][28] ),
    .A1(net2983),
    .S(net3209),
    .X(_00817_));
 sg13g2_mux2_1 _10723_ (.A0(\cpu.regs[11][29] ),
    .A1(net2982),
    .S(net3210),
    .X(_00818_));
 sg13g2_mux2_1 _10724_ (.A0(\cpu.regs[11][30] ),
    .A1(net3010),
    .S(net3210),
    .X(_00819_));
 sg13g2_mux2_1 _10725_ (.A0(\cpu.regs[11][31] ),
    .A1(net3008),
    .S(net3210),
    .X(_00820_));
 sg13g2_o21ai_1 _10726_ (.B1(net3701),
    .Y(_04910_),
    .A1(\cpu.Bimm[1] ),
    .A2(\cpu.Bimm[11] ));
 sg13g2_nand2_1 _10727_ (.Y(_04911_),
    .A(_04124_),
    .B(_04910_));
 sg13g2_nor2_1 _10728_ (.A(net3047),
    .B(net3203),
    .Y(_04912_));
 sg13g2_a21oi_1 _10729_ (.A1(_01687_),
    .A2(net3208),
    .Y(_00821_),
    .B1(_04912_));
 sg13g2_mux2_1 _10730_ (.A0(net3042),
    .A1(\cpu.regs[12][1] ),
    .S(net3208),
    .X(_00822_));
 sg13g2_mux2_1 _10731_ (.A0(net3039),
    .A1(\cpu.regs[12][2] ),
    .S(net3203),
    .X(_00823_));
 sg13g2_mux2_1 _10732_ (.A0(net3006),
    .A1(\cpu.regs[12][3] ),
    .S(net3205),
    .X(_00824_));
 sg13g2_mux2_1 _10733_ (.A0(net3004),
    .A1(\cpu.regs[12][4] ),
    .S(net3203),
    .X(_00825_));
 sg13g2_mux2_1 _10734_ (.A0(net3030),
    .A1(\cpu.regs[12][5] ),
    .S(net3206),
    .X(_00826_));
 sg13g2_mux2_1 _10735_ (.A0(net3038),
    .A1(\cpu.regs[12][6] ),
    .S(net3208),
    .X(_00827_));
 sg13g2_mux2_1 _10736_ (.A0(net3045),
    .A1(\cpu.regs[12][7] ),
    .S(net3205),
    .X(_00828_));
 sg13g2_mux2_1 _10737_ (.A0(net3028),
    .A1(\cpu.regs[12][8] ),
    .S(net3205),
    .X(_00829_));
 sg13g2_mux2_1 _10738_ (.A0(net3026),
    .A1(\cpu.regs[12][9] ),
    .S(net3205),
    .X(_00830_));
 sg13g2_mux2_1 _10739_ (.A0(net3024),
    .A1(\cpu.regs[12][10] ),
    .S(net3206),
    .X(_00831_));
 sg13g2_mux2_1 _10740_ (.A0(net3022),
    .A1(\cpu.regs[12][11] ),
    .S(net3206),
    .X(_00832_));
 sg13g2_mux2_1 _10741_ (.A0(net3001),
    .A1(\cpu.regs[12][12] ),
    .S(net3203),
    .X(_00833_));
 sg13g2_mux2_1 _10742_ (.A0(net3020),
    .A1(\cpu.regs[12][13] ),
    .S(net3203),
    .X(_00834_));
 sg13g2_nand2_1 _10743_ (.Y(_04913_),
    .A(\cpu.regs[12][14] ),
    .B(net3205));
 sg13g2_o21ai_1 _10744_ (.B1(_04913_),
    .Y(_00835_),
    .A1(net3036),
    .A2(net3205));
 sg13g2_nand2_1 _10745_ (.Y(_04914_),
    .A(\cpu.regs[12][15] ),
    .B(net3205));
 sg13g2_o21ai_1 _10746_ (.B1(_04914_),
    .Y(_00836_),
    .A1(net3034),
    .A2(net3205));
 sg13g2_mux2_1 _10747_ (.A0(net3000),
    .A1(\cpu.regs[12][16] ),
    .S(net3203),
    .X(_00837_));
 sg13g2_nand2_1 _10748_ (.Y(_04915_),
    .A(\cpu.regs[12][17] ),
    .B(net3206));
 sg13g2_o21ai_1 _10749_ (.B1(_04915_),
    .Y(_00838_),
    .A1(net2998),
    .A2(net3206));
 sg13g2_mux2_1 _10750_ (.A0(net2996),
    .A1(\cpu.regs[12][18] ),
    .S(net3207),
    .X(_00839_));
 sg13g2_nand2_1 _10751_ (.Y(_04916_),
    .A(\cpu.regs[12][19] ),
    .B(net3206));
 sg13g2_o21ai_1 _10752_ (.B1(_04916_),
    .Y(_00840_),
    .A1(net2994),
    .A2(net3206));
 sg13g2_mux2_1 _10753_ (.A0(net2991),
    .A1(\cpu.regs[12][20] ),
    .S(net3203),
    .X(_00841_));
 sg13g2_mux2_1 _10754_ (.A0(net2990),
    .A1(\cpu.regs[12][21] ),
    .S(net3207),
    .X(_00842_));
 sg13g2_mux2_1 _10755_ (.A0(net3017),
    .A1(\cpu.regs[12][22] ),
    .S(net3204),
    .X(_00843_));
 sg13g2_mux2_1 _10756_ (.A0(net3016),
    .A1(\cpu.regs[12][23] ),
    .S(net3204),
    .X(_00844_));
 sg13g2_mux2_1 _10757_ (.A0(net2987),
    .A1(\cpu.regs[12][24] ),
    .S(net3204),
    .X(_00845_));
 sg13g2_mux2_1 _10758_ (.A0(net2986),
    .A1(\cpu.regs[12][25] ),
    .S(net3207),
    .X(_00846_));
 sg13g2_mux2_1 _10759_ (.A0(net3014),
    .A1(\cpu.regs[12][26] ),
    .S(net3204),
    .X(_00847_));
 sg13g2_mux2_1 _10760_ (.A0(net3012),
    .A1(\cpu.regs[12][27] ),
    .S(net3204),
    .X(_00848_));
 sg13g2_mux2_1 _10761_ (.A0(net2983),
    .A1(\cpu.regs[12][28] ),
    .S(net3204),
    .X(_00849_));
 sg13g2_mux2_1 _10762_ (.A0(net2982),
    .A1(\cpu.regs[12][29] ),
    .S(net3204),
    .X(_00850_));
 sg13g2_mux2_1 _10763_ (.A0(net3010),
    .A1(\cpu.regs[12][30] ),
    .S(net3203),
    .X(_00851_));
 sg13g2_mux2_1 _10764_ (.A0(net3008),
    .A1(\cpu.regs[12][31] ),
    .S(net3204),
    .X(_00852_));
 sg13g2_nor3_2 _10765_ (.A(\cpu.Bimm[3] ),
    .B(_04122_),
    .C(_04895_),
    .Y(_04917_));
 sg13g2_nor2b_2 _10766_ (.A(_04903_),
    .B_N(_04917_),
    .Y(_04918_));
 sg13g2_mux2_1 _10767_ (.A0(\cpu.regs[7][0] ),
    .A1(net3046),
    .S(net3198),
    .X(_00853_));
 sg13g2_mux2_1 _10768_ (.A0(\cpu.regs[7][1] ),
    .A1(net3041),
    .S(net3198),
    .X(_00854_));
 sg13g2_mux2_1 _10769_ (.A0(\cpu.regs[7][2] ),
    .A1(net3040),
    .S(net3198),
    .X(_00855_));
 sg13g2_mux2_1 _10770_ (.A0(\cpu.regs[7][3] ),
    .A1(net3005),
    .S(net3200),
    .X(_00856_));
 sg13g2_mux2_1 _10771_ (.A0(\cpu.regs[7][4] ),
    .A1(net3003),
    .S(net3197),
    .X(_00857_));
 sg13g2_mux2_1 _10772_ (.A0(\cpu.regs[7][5] ),
    .A1(net3029),
    .S(net3201),
    .X(_00858_));
 sg13g2_mux2_1 _10773_ (.A0(\cpu.regs[7][6] ),
    .A1(net3037),
    .S(net3198),
    .X(_00859_));
 sg13g2_mux2_1 _10774_ (.A0(\cpu.regs[7][7] ),
    .A1(net3044),
    .S(net3200),
    .X(_00860_));
 sg13g2_mux2_1 _10775_ (.A0(\cpu.regs[7][8] ),
    .A1(net3027),
    .S(net3200),
    .X(_00861_));
 sg13g2_mux2_1 _10776_ (.A0(\cpu.regs[7][9] ),
    .A1(net3026),
    .S(net3200),
    .X(_00862_));
 sg13g2_mux2_1 _10777_ (.A0(\cpu.regs[7][10] ),
    .A1(net3023),
    .S(net3201),
    .X(_00863_));
 sg13g2_mux2_1 _10778_ (.A0(\cpu.regs[7][11] ),
    .A1(net3021),
    .S(net3201),
    .X(_00864_));
 sg13g2_mux2_1 _10779_ (.A0(\cpu.regs[7][12] ),
    .A1(net3002),
    .S(net3197),
    .X(_00865_));
 sg13g2_mux2_1 _10780_ (.A0(\cpu.regs[7][13] ),
    .A1(net3019),
    .S(net3197),
    .X(_00866_));
 sg13g2_nor2_1 _10781_ (.A(\cpu.regs[7][14] ),
    .B(net3200),
    .Y(_04919_));
 sg13g2_a21oi_1 _10782_ (.A1(net3035),
    .A2(net3200),
    .Y(_00867_),
    .B1(_04919_));
 sg13g2_nor2_1 _10783_ (.A(\cpu.regs[7][15] ),
    .B(net3200),
    .Y(_04920_));
 sg13g2_a21oi_1 _10784_ (.A1(net3033),
    .A2(net3200),
    .Y(_00868_),
    .B1(_04920_));
 sg13g2_mux2_1 _10785_ (.A0(\cpu.regs[7][16] ),
    .A1(net2999),
    .S(net3197),
    .X(_00869_));
 sg13g2_nor2_1 _10786_ (.A(\cpu.regs[7][17] ),
    .B(net3201),
    .Y(_04921_));
 sg13g2_a21oi_1 _10787_ (.A1(net2997),
    .A2(net3201),
    .Y(_00870_),
    .B1(_04921_));
 sg13g2_mux2_1 _10788_ (.A0(\cpu.regs[7][18] ),
    .A1(net2995),
    .S(net3199),
    .X(_00871_));
 sg13g2_nor2_1 _10789_ (.A(\cpu.regs[7][19] ),
    .B(net3199),
    .Y(_04922_));
 sg13g2_a21oi_1 _10790_ (.A1(net2993),
    .A2(net3199),
    .Y(_00872_),
    .B1(_04922_));
 sg13g2_mux2_1 _10791_ (.A0(\cpu.regs[7][20] ),
    .A1(net2992),
    .S(net3197),
    .X(_00873_));
 sg13g2_mux2_1 _10792_ (.A0(\cpu.regs[7][21] ),
    .A1(net2989),
    .S(net3202),
    .X(_00874_));
 sg13g2_mux2_1 _10793_ (.A0(\cpu.regs[7][22] ),
    .A1(net3018),
    .S(net3199),
    .X(_00875_));
 sg13g2_mux2_1 _10794_ (.A0(\cpu.regs[7][23] ),
    .A1(net3015),
    .S(net3202),
    .X(_00876_));
 sg13g2_mux2_1 _10795_ (.A0(\cpu.regs[7][24] ),
    .A1(net2988),
    .S(net3199),
    .X(_00877_));
 sg13g2_mux2_1 _10796_ (.A0(\cpu.regs[7][25] ),
    .A1(net2985),
    .S(net3202),
    .X(_00878_));
 sg13g2_mux2_1 _10797_ (.A0(\cpu.regs[7][26] ),
    .A1(net3013),
    .S(net3197),
    .X(_00879_));
 sg13g2_mux2_1 _10798_ (.A0(\cpu.regs[7][27] ),
    .A1(net3011),
    .S(net3199),
    .X(_00880_));
 sg13g2_mux2_1 _10799_ (.A0(\cpu.regs[7][28] ),
    .A1(net2984),
    .S(net3199),
    .X(_00881_));
 sg13g2_mux2_1 _10800_ (.A0(\cpu.regs[7][29] ),
    .A1(net2981),
    .S(net3199),
    .X(_00882_));
 sg13g2_mux2_1 _10801_ (.A0(\cpu.regs[7][30] ),
    .A1(net3009),
    .S(net3197),
    .X(_00883_));
 sg13g2_mux2_1 _10802_ (.A0(\cpu.regs[7][31] ),
    .A1(net3007),
    .S(net3197),
    .X(_00884_));
 sg13g2_and3_1 _10803_ (.X(_04923_),
    .A(\cpu.Bimm[1] ),
    .B(_01690_),
    .C(net3701));
 sg13g2_nand2_2 _10804_ (.Y(_04924_),
    .A(_04897_),
    .B(_04923_));
 sg13g2_mux2_1 _10805_ (.A0(net3046),
    .A1(\cpu.regs[2][0] ),
    .S(net3196),
    .X(_00885_));
 sg13g2_mux2_1 _10806_ (.A0(net3041),
    .A1(\cpu.regs[2][1] ),
    .S(net3196),
    .X(_00886_));
 sg13g2_mux2_1 _10807_ (.A0(net3040),
    .A1(\cpu.regs[2][2] ),
    .S(net3196),
    .X(_00887_));
 sg13g2_mux2_1 _10808_ (.A0(net3005),
    .A1(\cpu.regs[2][3] ),
    .S(net3195),
    .X(_00888_));
 sg13g2_mux2_1 _10809_ (.A0(net3003),
    .A1(\cpu.regs[2][4] ),
    .S(net3196),
    .X(_00889_));
 sg13g2_mux2_1 _10810_ (.A0(net3029),
    .A1(\cpu.regs[2][5] ),
    .S(net3195),
    .X(_00890_));
 sg13g2_mux2_1 _10811_ (.A0(net3038),
    .A1(\cpu.regs[2][6] ),
    .S(net3196),
    .X(_00891_));
 sg13g2_mux2_1 _10812_ (.A0(net3044),
    .A1(\cpu.regs[2][7] ),
    .S(net3194),
    .X(_00892_));
 sg13g2_mux2_1 _10813_ (.A0(net3027),
    .A1(\cpu.regs[2][8] ),
    .S(net3195),
    .X(_00893_));
 sg13g2_mux2_1 _10814_ (.A0(net3025),
    .A1(\cpu.regs[2][9] ),
    .S(net3195),
    .X(_00894_));
 sg13g2_mux2_1 _10815_ (.A0(net3023),
    .A1(\cpu.regs[2][10] ),
    .S(net3195),
    .X(_00895_));
 sg13g2_mux2_1 _10816_ (.A0(net3021),
    .A1(\cpu.regs[2][11] ),
    .S(net3194),
    .X(_00896_));
 sg13g2_mux2_1 _10817_ (.A0(net3001),
    .A1(\cpu.regs[2][12] ),
    .S(net3193),
    .X(_00897_));
 sg13g2_mux2_1 _10818_ (.A0(net3019),
    .A1(\cpu.regs[2][13] ),
    .S(net3193),
    .X(_00898_));
 sg13g2_nand2_1 _10819_ (.Y(_04925_),
    .A(\cpu.regs[2][14] ),
    .B(net3194));
 sg13g2_o21ai_1 _10820_ (.B1(_04925_),
    .Y(_00899_),
    .A1(net3035),
    .A2(net3194));
 sg13g2_nand2_1 _10821_ (.Y(_04926_),
    .A(\cpu.regs[2][15] ),
    .B(net3194));
 sg13g2_o21ai_1 _10822_ (.B1(_04926_),
    .Y(_00900_),
    .A1(net3033),
    .A2(net3194));
 sg13g2_mux2_1 _10823_ (.A0(net2999),
    .A1(\cpu.regs[2][16] ),
    .S(net3196),
    .X(_00901_));
 sg13g2_nand2_1 _10824_ (.Y(_04927_),
    .A(\cpu.regs[2][17] ),
    .B(net3194));
 sg13g2_o21ai_1 _10825_ (.B1(_04927_),
    .Y(_00902_),
    .A1(net2997),
    .A2(net3194));
 sg13g2_mux2_1 _10826_ (.A0(net2995),
    .A1(\cpu.regs[2][18] ),
    .S(net3191),
    .X(_00903_));
 sg13g2_nand2_1 _10827_ (.Y(_04928_),
    .A(\cpu.regs[2][19] ),
    .B(net3191));
 sg13g2_o21ai_1 _10828_ (.B1(_04928_),
    .Y(_00904_),
    .A1(net2993),
    .A2(net3191));
 sg13g2_mux2_1 _10829_ (.A0(net2991),
    .A1(\cpu.regs[2][20] ),
    .S(net3193),
    .X(_00905_));
 sg13g2_mux2_1 _10830_ (.A0(net2989),
    .A1(\cpu.regs[2][21] ),
    .S(net3192),
    .X(_00906_));
 sg13g2_mux2_1 _10831_ (.A0(net3018),
    .A1(\cpu.regs[2][22] ),
    .S(net3191),
    .X(_00907_));
 sg13g2_mux2_1 _10832_ (.A0(net3015),
    .A1(\cpu.regs[2][23] ),
    .S(net3192),
    .X(_00908_));
 sg13g2_mux2_1 _10833_ (.A0(net2988),
    .A1(\cpu.regs[2][24] ),
    .S(net3191),
    .X(_00909_));
 sg13g2_mux2_1 _10834_ (.A0(net2985),
    .A1(\cpu.regs[2][25] ),
    .S(net3191),
    .X(_00910_));
 sg13g2_mux2_1 _10835_ (.A0(net3013),
    .A1(\cpu.regs[2][26] ),
    .S(net3193),
    .X(_00911_));
 sg13g2_mux2_1 _10836_ (.A0(net3011),
    .A1(\cpu.regs[2][27] ),
    .S(net3192),
    .X(_00912_));
 sg13g2_mux2_1 _10837_ (.A0(net2984),
    .A1(\cpu.regs[2][28] ),
    .S(net3191),
    .X(_00913_));
 sg13g2_mux2_1 _10838_ (.A0(net2981),
    .A1(\cpu.regs[2][29] ),
    .S(net3191),
    .X(_00914_));
 sg13g2_mux2_1 _10839_ (.A0(net3009),
    .A1(\cpu.regs[2][30] ),
    .S(net3193),
    .X(_00915_));
 sg13g2_mux2_1 _10840_ (.A0(net3007),
    .A1(\cpu.regs[2][31] ),
    .S(net3193),
    .X(_00916_));
 sg13g2_nor3_2 _10841_ (.A(_02579_),
    .B(_03452_),
    .C(_04867_),
    .Y(_04929_));
 sg13g2_mux2_1 _10842_ (.A0(\irqvect[0][0] ),
    .A1(net3326),
    .S(net3074),
    .X(_00917_));
 sg13g2_mux2_1 _10843_ (.A0(\irqvect[0][1] ),
    .A1(net3327),
    .S(net3076),
    .X(_00918_));
 sg13g2_nor2_1 _10844_ (.A(\irqvect[0][2] ),
    .B(net3075),
    .Y(_04930_));
 sg13g2_a21oi_1 _10845_ (.A1(_02928_),
    .A2(net3074),
    .Y(_00919_),
    .B1(_04930_));
 sg13g2_mux2_1 _10846_ (.A0(\irqvect[0][3] ),
    .A1(net3328),
    .S(net3076),
    .X(_00920_));
 sg13g2_mux2_1 _10847_ (.A0(\irqvect[0][4] ),
    .A1(net3329),
    .S(net3075),
    .X(_00921_));
 sg13g2_mux2_1 _10848_ (.A0(\irqvect[0][5] ),
    .A1(net3330),
    .S(net3075),
    .X(_00922_));
 sg13g2_nor2_1 _10849_ (.A(\irqvect[0][6] ),
    .B(net3075),
    .Y(_04931_));
 sg13g2_a21oi_1 _10850_ (.A1(_03267_),
    .A2(net3075),
    .Y(_00923_),
    .B1(_04931_));
 sg13g2_nor2_1 _10851_ (.A(\irqvect[0][7] ),
    .B(net3075),
    .Y(_04932_));
 sg13g2_a21oi_1 _10852_ (.A1(_03193_),
    .A2(net3075),
    .Y(_00924_),
    .B1(_04932_));
 sg13g2_nor2_1 _10853_ (.A(\irqvect[0][8] ),
    .B(net3077),
    .Y(_04933_));
 sg13g2_a21oi_1 _10854_ (.A1(_03120_),
    .A2(net3076),
    .Y(_00925_),
    .B1(_04933_));
 sg13g2_nor2_1 _10855_ (.A(\irqvect[0][9] ),
    .B(net3077),
    .Y(_04934_));
 sg13g2_a21oi_1 _10856_ (.A1(_03033_),
    .A2(net3077),
    .Y(_00926_),
    .B1(_04934_));
 sg13g2_nor2_1 _10857_ (.A(\irqvect[0][10] ),
    .B(net3076),
    .Y(_04935_));
 sg13g2_a21oi_1 _10858_ (.A1(_02947_),
    .A2(net3076),
    .Y(_00927_),
    .B1(_04935_));
 sg13g2_nor2_1 _10859_ (.A(\irqvect[0][11] ),
    .B(net3073),
    .Y(_04936_));
 sg13g2_a21oi_1 _10860_ (.A1(_02861_),
    .A2(net3073),
    .Y(_00928_),
    .B1(_04936_));
 sg13g2_nor2_1 _10861_ (.A(\irqvect[0][12] ),
    .B(net3072),
    .Y(_04937_));
 sg13g2_a21oi_1 _10862_ (.A1(_02778_),
    .A2(net3072),
    .Y(_00929_),
    .B1(_04937_));
 sg13g2_nor2_1 _10863_ (.A(\irqvect[0][13] ),
    .B(net3077),
    .Y(_04938_));
 sg13g2_a21oi_1 _10864_ (.A1(_02682_),
    .A2(net3077),
    .Y(_00930_),
    .B1(_04938_));
 sg13g2_nor2_1 _10865_ (.A(\irqvect[0][14] ),
    .B(net3074),
    .Y(_04939_));
 sg13g2_a21oi_1 _10866_ (.A1(_03288_),
    .A2(net3074),
    .Y(_00931_),
    .B1(_04939_));
 sg13g2_nor2_1 _10867_ (.A(\irqvect[0][15] ),
    .B(net3074),
    .Y(_04940_));
 sg13g2_a21oi_1 _10868_ (.A1(_03216_),
    .A2(net3074),
    .Y(_00932_),
    .B1(_04940_));
 sg13g2_nor2_1 _10869_ (.A(\irqvect[0][16] ),
    .B(net3074),
    .Y(_04941_));
 sg13g2_a21oi_1 _10870_ (.A1(_03142_),
    .A2(net3074),
    .Y(_00933_),
    .B1(_04941_));
 sg13g2_nor2_1 _10871_ (.A(\irqvect[0][17] ),
    .B(net3071),
    .Y(_04942_));
 sg13g2_a21oi_1 _10872_ (.A1(_03054_),
    .A2(net3070),
    .Y(_00934_),
    .B1(_04942_));
 sg13g2_nor2_1 _10873_ (.A(\irqvect[0][18] ),
    .B(net3070),
    .Y(_04943_));
 sg13g2_a21oi_1 _10874_ (.A1(_02967_),
    .A2(net3070),
    .Y(_00935_),
    .B1(_04943_));
 sg13g2_nor2_1 _10875_ (.A(\irqvect[0][19] ),
    .B(net3073),
    .Y(_04944_));
 sg13g2_a21oi_1 _10876_ (.A1(_02881_),
    .A2(net3073),
    .Y(_00936_),
    .B1(_04944_));
 sg13g2_nor2_1 _10877_ (.A(\irqvect[0][20] ),
    .B(net3070),
    .Y(_04945_));
 sg13g2_a21oi_1 _10878_ (.A1(_02798_),
    .A2(net3070),
    .Y(_00937_),
    .B1(_04945_));
 sg13g2_nor2_1 _10879_ (.A(\irqvect[0][21] ),
    .B(net3072),
    .Y(_04946_));
 sg13g2_a21oi_1 _10880_ (.A1(_02703_),
    .A2(net3072),
    .Y(_00938_),
    .B1(_04946_));
 sg13g2_nor2_1 _10881_ (.A(\irqvect[0][22] ),
    .B(net3071),
    .Y(_04947_));
 sg13g2_a21oi_1 _10882_ (.A1(_03269_),
    .A2(net3070),
    .Y(_00939_),
    .B1(_04947_));
 sg13g2_nor2_1 _10883_ (.A(\irqvect[0][23] ),
    .B(net3071),
    .Y(_04948_));
 sg13g2_a21oi_1 _10884_ (.A1(_03195_),
    .A2(net3071),
    .Y(_00940_),
    .B1(_04948_));
 sg13g2_nor2_1 _10885_ (.A(\irqvect[0][24] ),
    .B(net3071),
    .Y(_04949_));
 sg13g2_a21oi_1 _10886_ (.A1(_03122_),
    .A2(net3071),
    .Y(_00941_),
    .B1(_04949_));
 sg13g2_nor2_1 _10887_ (.A(\irqvect[0][25] ),
    .B(net3076),
    .Y(_04950_));
 sg13g2_a21oi_1 _10888_ (.A1(_03035_),
    .A2(net3076),
    .Y(_00942_),
    .B1(_04950_));
 sg13g2_nor2_1 _10889_ (.A(\irqvect[0][26] ),
    .B(net3070),
    .Y(_04951_));
 sg13g2_a21oi_1 _10890_ (.A1(_02949_),
    .A2(net3070),
    .Y(_00943_),
    .B1(_04951_));
 sg13g2_nor2_1 _10891_ (.A(\irqvect[0][27] ),
    .B(net3072),
    .Y(_04952_));
 sg13g2_a21oi_1 _10892_ (.A1(_02863_),
    .A2(net3072),
    .Y(_00944_),
    .B1(_04952_));
 sg13g2_nor2_1 _10893_ (.A(\irqvect[0][28] ),
    .B(net3073),
    .Y(_04953_));
 sg13g2_a21oi_1 _10894_ (.A1(_02780_),
    .A2(net3073),
    .Y(_00945_),
    .B1(_04953_));
 sg13g2_nor2_1 _10895_ (.A(\irqvect[0][29] ),
    .B(net3073),
    .Y(_04954_));
 sg13g2_a21oi_1 _10896_ (.A1(_02684_),
    .A2(net3073),
    .Y(_00946_),
    .B1(_04954_));
 sg13g2_and2_1 _10897_ (.A(_04904_),
    .B(_04923_),
    .X(_04955_));
 sg13g2_mux2_1 _10898_ (.A0(\cpu.regs[10][0] ),
    .A1(net3047),
    .S(net3189),
    .X(_00947_));
 sg13g2_mux2_1 _10899_ (.A0(\cpu.regs[10][1] ),
    .A1(net3042),
    .S(net3189),
    .X(_00948_));
 sg13g2_mux2_1 _10900_ (.A0(\cpu.regs[10][2] ),
    .A1(net3039),
    .S(net3189),
    .X(_00949_));
 sg13g2_mux2_1 _10901_ (.A0(\cpu.regs[10][3] ),
    .A1(net3006),
    .S(net3188),
    .X(_00950_));
 sg13g2_mux2_1 _10902_ (.A0(\cpu.regs[10][4] ),
    .A1(net3004),
    .S(net3189),
    .X(_00951_));
 sg13g2_mux2_1 _10903_ (.A0(\cpu.regs[10][5] ),
    .A1(net3030),
    .S(net3188),
    .X(_00952_));
 sg13g2_mux2_1 _10904_ (.A0(\cpu.regs[10][6] ),
    .A1(net3038),
    .S(net3189),
    .X(_00953_));
 sg13g2_mux2_1 _10905_ (.A0(\cpu.regs[10][7] ),
    .A1(net3045),
    .S(net3188),
    .X(_00954_));
 sg13g2_mux2_1 _10906_ (.A0(\cpu.regs[10][8] ),
    .A1(net3028),
    .S(net3188),
    .X(_00955_));
 sg13g2_mux2_1 _10907_ (.A0(\cpu.regs[10][9] ),
    .A1(net3025),
    .S(net3189),
    .X(_00956_));
 sg13g2_mux2_1 _10908_ (.A0(\cpu.regs[10][10] ),
    .A1(net3024),
    .S(net3188),
    .X(_00957_));
 sg13g2_mux2_1 _10909_ (.A0(\cpu.regs[10][11] ),
    .A1(net3022),
    .S(net3187),
    .X(_00958_));
 sg13g2_mux2_1 _10910_ (.A0(\cpu.regs[10][12] ),
    .A1(net3002),
    .S(net3186),
    .X(_00959_));
 sg13g2_mux2_1 _10911_ (.A0(\cpu.regs[10][13] ),
    .A1(net3020),
    .S(net3186),
    .X(_00960_));
 sg13g2_nor2_1 _10912_ (.A(\cpu.regs[10][14] ),
    .B(net3187),
    .Y(_04956_));
 sg13g2_a21oi_1 _10913_ (.A1(net3036),
    .A2(net3187),
    .Y(_00961_),
    .B1(_04956_));
 sg13g2_nor2_1 _10914_ (.A(\cpu.regs[10][15] ),
    .B(net3187),
    .Y(_04957_));
 sg13g2_a21oi_1 _10915_ (.A1(net3034),
    .A2(net3187),
    .Y(_00962_),
    .B1(_04957_));
 sg13g2_mux2_1 _10916_ (.A0(\cpu.regs[10][16] ),
    .A1(net3000),
    .S(net3189),
    .X(_00963_));
 sg13g2_nor2_1 _10917_ (.A(\cpu.regs[10][17] ),
    .B(net3187),
    .Y(_04958_));
 sg13g2_a21oi_1 _10918_ (.A1(net2998),
    .A2(net3187),
    .Y(_00964_),
    .B1(_04958_));
 sg13g2_mux2_1 _10919_ (.A0(\cpu.regs[10][18] ),
    .A1(net2996),
    .S(net3187),
    .X(_00965_));
 sg13g2_nor2_1 _10920_ (.A(\cpu.regs[10][19] ),
    .B(net3185),
    .Y(_04959_));
 sg13g2_a21oi_1 _10921_ (.A1(net2994),
    .A2(net3185),
    .Y(_00966_),
    .B1(_04959_));
 sg13g2_mux2_1 _10922_ (.A0(\cpu.regs[10][20] ),
    .A1(net2992),
    .S(net3186),
    .X(_00967_));
 sg13g2_mux2_1 _10923_ (.A0(\cpu.regs[10][21] ),
    .A1(net2989),
    .S(net3185),
    .X(_00968_));
 sg13g2_mux2_1 _10924_ (.A0(\cpu.regs[10][22] ),
    .A1(net3017),
    .S(net3185),
    .X(_00969_));
 sg13g2_mux2_1 _10925_ (.A0(\cpu.regs[10][23] ),
    .A1(net3016),
    .S(net3185),
    .X(_00970_));
 sg13g2_mux2_1 _10926_ (.A0(\cpu.regs[10][24] ),
    .A1(net2987),
    .S(net3185),
    .X(_00971_));
 sg13g2_mux2_1 _10927_ (.A0(\cpu.regs[10][25] ),
    .A1(net2986),
    .S(net3185),
    .X(_00972_));
 sg13g2_mux2_1 _10928_ (.A0(\cpu.regs[10][26] ),
    .A1(net3014),
    .S(net3186),
    .X(_00973_));
 sg13g2_mux2_1 _10929_ (.A0(\cpu.regs[10][27] ),
    .A1(net3012),
    .S(net3185),
    .X(_00974_));
 sg13g2_mux2_1 _10930_ (.A0(\cpu.regs[10][28] ),
    .A1(net2983),
    .S(net3186),
    .X(_00975_));
 sg13g2_mux2_1 _10931_ (.A0(\cpu.regs[10][29] ),
    .A1(net2982),
    .S(net3190),
    .X(_00976_));
 sg13g2_mux2_1 _10932_ (.A0(\cpu.regs[10][30] ),
    .A1(net3010),
    .S(net3186),
    .X(_00977_));
 sg13g2_mux2_1 _10933_ (.A0(\cpu.regs[10][31] ),
    .A1(net3008),
    .S(net3186),
    .X(_00978_));
 sg13g2_nor3_2 _10934_ (.A(net3125),
    .B(_03443_),
    .C(_04868_),
    .Y(_04960_));
 sg13g2_mux2_1 _10935_ (.A0(\irqvect[2][0] ),
    .A1(net3326),
    .S(net3067),
    .X(_00979_));
 sg13g2_mux2_1 _10936_ (.A0(\irqvect[2][1] ),
    .A1(net3327),
    .S(net3068),
    .X(_00980_));
 sg13g2_nor2_1 _10937_ (.A(\irqvect[2][2] ),
    .B(net3067),
    .Y(_04961_));
 sg13g2_a21oi_1 _10938_ (.A1(_02928_),
    .A2(net3067),
    .Y(_00981_),
    .B1(_04961_));
 sg13g2_mux2_1 _10939_ (.A0(\irqvect[2][3] ),
    .A1(net3328),
    .S(net3068),
    .X(_00982_));
 sg13g2_mux2_1 _10940_ (.A0(\irqvect[2][4] ),
    .A1(net3329),
    .S(net3068),
    .X(_00983_));
 sg13g2_mux2_1 _10941_ (.A0(\irqvect[2][5] ),
    .A1(net3330),
    .S(net3068),
    .X(_00984_));
 sg13g2_nor2_1 _10942_ (.A(\irqvect[2][6] ),
    .B(net3068),
    .Y(_04962_));
 sg13g2_a21oi_1 _10943_ (.A1(_03267_),
    .A2(net3068),
    .Y(_00985_),
    .B1(_04962_));
 sg13g2_nor2_1 _10944_ (.A(\irqvect[2][7] ),
    .B(net3067),
    .Y(_04963_));
 sg13g2_a21oi_1 _10945_ (.A1(_03193_),
    .A2(net3068),
    .Y(_00986_),
    .B1(_04963_));
 sg13g2_nor2_1 _10946_ (.A(\irqvect[2][8] ),
    .B(net3069),
    .Y(_04964_));
 sg13g2_a21oi_1 _10947_ (.A1(_03120_),
    .A2(net3069),
    .Y(_00987_),
    .B1(_04964_));
 sg13g2_nor2_1 _10948_ (.A(\irqvect[2][9] ),
    .B(net3066),
    .Y(_04965_));
 sg13g2_a21oi_1 _10949_ (.A1(_03033_),
    .A2(net3064),
    .Y(_00988_),
    .B1(_04965_));
 sg13g2_nor2_1 _10950_ (.A(\irqvect[2][10] ),
    .B(net3067),
    .Y(_04966_));
 sg13g2_a21oi_1 _10951_ (.A1(_02947_),
    .A2(net3067),
    .Y(_00989_),
    .B1(_04966_));
 sg13g2_nor2_1 _10952_ (.A(\irqvect[2][11] ),
    .B(net3062),
    .Y(_04967_));
 sg13g2_a21oi_1 _10953_ (.A1(_02861_),
    .A2(net3062),
    .Y(_00990_),
    .B1(_04967_));
 sg13g2_nor2_1 _10954_ (.A(\irqvect[2][12] ),
    .B(net3066),
    .Y(_04968_));
 sg13g2_a21oi_1 _10955_ (.A1(_02778_),
    .A2(net3066),
    .Y(_00991_),
    .B1(_04968_));
 sg13g2_nor2_1 _10956_ (.A(\irqvect[2][13] ),
    .B(net3069),
    .Y(_04969_));
 sg13g2_a21oi_1 _10957_ (.A1(_02682_),
    .A2(net3069),
    .Y(_00992_),
    .B1(_04969_));
 sg13g2_nor2_1 _10958_ (.A(\irqvect[2][14] ),
    .B(net3067),
    .Y(_04970_));
 sg13g2_a21oi_1 _10959_ (.A1(_03288_),
    .A2(net3067),
    .Y(_00993_),
    .B1(_04970_));
 sg13g2_nor2_1 _10960_ (.A(\irqvect[2][15] ),
    .B(net3062),
    .Y(_04971_));
 sg13g2_a21oi_1 _10961_ (.A1(_03216_),
    .A2(net3062),
    .Y(_00994_),
    .B1(_04971_));
 sg13g2_nor2_1 _10962_ (.A(\irqvect[2][16] ),
    .B(net3062),
    .Y(_04972_));
 sg13g2_a21oi_1 _10963_ (.A1(_03142_),
    .A2(net3062),
    .Y(_00995_),
    .B1(_04972_));
 sg13g2_nor2_1 _10964_ (.A(\irqvect[2][17] ),
    .B(net3065),
    .Y(_04973_));
 sg13g2_a21oi_1 _10965_ (.A1(_03054_),
    .A2(net3065),
    .Y(_00996_),
    .B1(_04973_));
 sg13g2_nor2_1 _10966_ (.A(\irqvect[2][18] ),
    .B(net3065),
    .Y(_04974_));
 sg13g2_a21oi_1 _10967_ (.A1(_02967_),
    .A2(net3065),
    .Y(_00997_),
    .B1(_04974_));
 sg13g2_nor2_1 _10968_ (.A(\irqvect[2][19] ),
    .B(net3063),
    .Y(_04975_));
 sg13g2_a21oi_1 _10969_ (.A1(_02881_),
    .A2(net3063),
    .Y(_00998_),
    .B1(_04975_));
 sg13g2_nor2_1 _10970_ (.A(\irqvect[2][20] ),
    .B(net3065),
    .Y(_04976_));
 sg13g2_a21oi_1 _10971_ (.A1(_02798_),
    .A2(net3065),
    .Y(_00999_),
    .B1(_04976_));
 sg13g2_nor2_1 _10972_ (.A(\irqvect[2][21] ),
    .B(net3066),
    .Y(_04977_));
 sg13g2_a21oi_1 _10973_ (.A1(_02703_),
    .A2(net3066),
    .Y(_01000_),
    .B1(_04977_));
 sg13g2_nor2_1 _10974_ (.A(\irqvect[2][22] ),
    .B(net3064),
    .Y(_04978_));
 sg13g2_a21oi_1 _10975_ (.A1(_03269_),
    .A2(net3064),
    .Y(_01001_),
    .B1(_04978_));
 sg13g2_nor2_1 _10976_ (.A(\irqvect[2][23] ),
    .B(net3064),
    .Y(_04979_));
 sg13g2_a21oi_1 _10977_ (.A1(_03195_),
    .A2(net3064),
    .Y(_01002_),
    .B1(_04979_));
 sg13g2_nor2_1 _10978_ (.A(\irqvect[2][24] ),
    .B(net3064),
    .Y(_04980_));
 sg13g2_a21oi_1 _10979_ (.A1(_03122_),
    .A2(net3064),
    .Y(_01003_),
    .B1(_04980_));
 sg13g2_nor2_1 _10980_ (.A(\irqvect[2][25] ),
    .B(net3069),
    .Y(_04981_));
 sg13g2_a21oi_1 _10981_ (.A1(_03035_),
    .A2(net3069),
    .Y(_01004_),
    .B1(_04981_));
 sg13g2_nor2_1 _10982_ (.A(\irqvect[2][26] ),
    .B(net3064),
    .Y(_04982_));
 sg13g2_a21oi_1 _10983_ (.A1(_02949_),
    .A2(net3065),
    .Y(_01005_),
    .B1(_04982_));
 sg13g2_nor2_1 _10984_ (.A(\irqvect[2][27] ),
    .B(net3066),
    .Y(_04983_));
 sg13g2_a21oi_1 _10985_ (.A1(_02863_),
    .A2(net3066),
    .Y(_01006_),
    .B1(_04983_));
 sg13g2_nor2_1 _10986_ (.A(\irqvect[2][28] ),
    .B(net3062),
    .Y(_04984_));
 sg13g2_a21oi_1 _10987_ (.A1(_02780_),
    .A2(net3062),
    .Y(_01007_),
    .B1(_04984_));
 sg13g2_nor2_1 _10988_ (.A(\irqvect[2][29] ),
    .B(net3063),
    .Y(_04985_));
 sg13g2_a21oi_1 _10989_ (.A1(_02684_),
    .A2(net3063),
    .Y(_01008_),
    .B1(_04985_));
 sg13g2_nand2_1 _10990_ (.Y(_04986_),
    .A(_04124_),
    .B(_04923_));
 sg13g2_nor2_1 _10991_ (.A(net3047),
    .B(net3184),
    .Y(_04987_));
 sg13g2_a21oi_1 _10992_ (.A1(_01688_),
    .A2(net3184),
    .Y(_01009_),
    .B1(_04987_));
 sg13g2_mux2_1 _10993_ (.A0(net3042),
    .A1(\cpu.regs[14][1] ),
    .S(net3184),
    .X(_01010_));
 sg13g2_mux2_1 _10994_ (.A0(net3039),
    .A1(\cpu.regs[14][2] ),
    .S(net3179),
    .X(_01011_));
 sg13g2_mux2_1 _10995_ (.A0(net3006),
    .A1(\cpu.regs[14][3] ),
    .S(net3182),
    .X(_01012_));
 sg13g2_mux2_1 _10996_ (.A0(net3004),
    .A1(\cpu.regs[14][4] ),
    .S(net3179),
    .X(_01013_));
 sg13g2_mux2_1 _10997_ (.A0(net3030),
    .A1(\cpu.regs[14][5] ),
    .S(net3183),
    .X(_01014_));
 sg13g2_mux2_1 _10998_ (.A0(net3038),
    .A1(\cpu.regs[14][6] ),
    .S(net3179),
    .X(_01015_));
 sg13g2_mux2_1 _10999_ (.A0(net3045),
    .A1(\cpu.regs[14][7] ),
    .S(net3182),
    .X(_01016_));
 sg13g2_mux2_1 _11000_ (.A0(net3028),
    .A1(\cpu.regs[14][8] ),
    .S(net3182),
    .X(_01017_));
 sg13g2_mux2_1 _11001_ (.A0(net3025),
    .A1(\cpu.regs[14][9] ),
    .S(net3182),
    .X(_01018_));
 sg13g2_mux2_1 _11002_ (.A0(net3024),
    .A1(\cpu.regs[14][10] ),
    .S(net3183),
    .X(_01019_));
 sg13g2_mux2_1 _11003_ (.A0(net3022),
    .A1(\cpu.regs[14][11] ),
    .S(net3183),
    .X(_01020_));
 sg13g2_mux2_1 _11004_ (.A0(net3001),
    .A1(\cpu.regs[14][12] ),
    .S(net3179),
    .X(_01021_));
 sg13g2_mux2_1 _11005_ (.A0(net3020),
    .A1(\cpu.regs[14][13] ),
    .S(net3179),
    .X(_01022_));
 sg13g2_nand2_1 _11006_ (.Y(_04988_),
    .A(\cpu.regs[14][14] ),
    .B(net3183));
 sg13g2_o21ai_1 _11007_ (.B1(_04988_),
    .Y(_01023_),
    .A1(net3036),
    .A2(net3182));
 sg13g2_nand2_1 _11008_ (.Y(_04989_),
    .A(\cpu.regs[14][15] ),
    .B(net3182));
 sg13g2_o21ai_1 _11009_ (.B1(_04989_),
    .Y(_01024_),
    .A1(net3034),
    .A2(net3182));
 sg13g2_mux2_1 _11010_ (.A0(net3000),
    .A1(\cpu.regs[14][16] ),
    .S(net3179),
    .X(_01025_));
 sg13g2_nand2_1 _11011_ (.Y(_04990_),
    .A(\cpu.regs[14][17] ),
    .B(net3183));
 sg13g2_o21ai_1 _11012_ (.B1(_04990_),
    .Y(_01026_),
    .A1(net2998),
    .A2(net3183));
 sg13g2_mux2_1 _11013_ (.A0(net2996),
    .A1(\cpu.regs[14][18] ),
    .S(net3181),
    .X(_01027_));
 sg13g2_nand2_1 _11014_ (.Y(_04991_),
    .A(\cpu.regs[14][19] ),
    .B(net3180));
 sg13g2_o21ai_1 _11015_ (.B1(_04991_),
    .Y(_01028_),
    .A1(net2994),
    .A2(net3180));
 sg13g2_mux2_1 _11016_ (.A0(net2991),
    .A1(\cpu.regs[14][20] ),
    .S(net3179),
    .X(_01029_));
 sg13g2_mux2_1 _11017_ (.A0(net2990),
    .A1(\cpu.regs[14][21] ),
    .S(net3181),
    .X(_01030_));
 sg13g2_mux2_1 _11018_ (.A0(net3017),
    .A1(\cpu.regs[14][22] ),
    .S(net3180),
    .X(_01031_));
 sg13g2_mux2_1 _11019_ (.A0(net3015),
    .A1(\cpu.regs[14][23] ),
    .S(net3181),
    .X(_01032_));
 sg13g2_mux2_1 _11020_ (.A0(net2987),
    .A1(\cpu.regs[14][24] ),
    .S(net3180),
    .X(_01033_));
 sg13g2_mux2_1 _11021_ (.A0(net2986),
    .A1(\cpu.regs[14][25] ),
    .S(net3181),
    .X(_01034_));
 sg13g2_mux2_1 _11022_ (.A0(net3014),
    .A1(\cpu.regs[14][26] ),
    .S(net3180),
    .X(_01035_));
 sg13g2_mux2_1 _11023_ (.A0(net3011),
    .A1(\cpu.regs[14][27] ),
    .S(net3180),
    .X(_01036_));
 sg13g2_mux2_1 _11024_ (.A0(net2983),
    .A1(\cpu.regs[14][28] ),
    .S(net3180),
    .X(_01037_));
 sg13g2_mux2_1 _11025_ (.A0(net2982),
    .A1(\cpu.regs[14][29] ),
    .S(net3182),
    .X(_01038_));
 sg13g2_mux2_1 _11026_ (.A0(net3010),
    .A1(\cpu.regs[14][30] ),
    .S(net3179),
    .X(_01039_));
 sg13g2_mux2_1 _11027_ (.A0(net3008),
    .A1(\cpu.regs[14][31] ),
    .S(net3180),
    .X(_01040_));
 sg13g2_and2_1 _11028_ (.A(_04917_),
    .B(_04923_),
    .X(_04992_));
 sg13g2_mux2_1 _11029_ (.A0(\cpu.regs[6][0] ),
    .A1(net3046),
    .S(net3174),
    .X(_01041_));
 sg13g2_mux2_1 _11030_ (.A0(\cpu.regs[6][1] ),
    .A1(net3041),
    .S(net3174),
    .X(_01042_));
 sg13g2_mux2_1 _11031_ (.A0(\cpu.regs[6][2] ),
    .A1(net3040),
    .S(net3173),
    .X(_01043_));
 sg13g2_mux2_1 _11032_ (.A0(\cpu.regs[6][3] ),
    .A1(net3005),
    .S(net3177),
    .X(_01044_));
 sg13g2_mux2_1 _11033_ (.A0(\cpu.regs[6][4] ),
    .A1(net3003),
    .S(net3174),
    .X(_01045_));
 sg13g2_mux2_1 _11034_ (.A0(\cpu.regs[6][5] ),
    .A1(net3029),
    .S(net3176),
    .X(_01046_));
 sg13g2_mux2_1 _11035_ (.A0(\cpu.regs[6][6] ),
    .A1(net3037),
    .S(net3174),
    .X(_01047_));
 sg13g2_mux2_1 _11036_ (.A0(\cpu.regs[6][7] ),
    .A1(net3044),
    .S(net3176),
    .X(_01048_));
 sg13g2_mux2_1 _11037_ (.A0(\cpu.regs[6][8] ),
    .A1(net3027),
    .S(net3176),
    .X(_01049_));
 sg13g2_mux2_1 _11038_ (.A0(\cpu.regs[6][9] ),
    .A1(net3026),
    .S(net3176),
    .X(_01050_));
 sg13g2_mux2_1 _11039_ (.A0(\cpu.regs[6][10] ),
    .A1(net3023),
    .S(net3177),
    .X(_01051_));
 sg13g2_mux2_1 _11040_ (.A0(\cpu.regs[6][11] ),
    .A1(net3021),
    .S(net3177),
    .X(_01052_));
 sg13g2_mux2_1 _11041_ (.A0(\cpu.regs[6][12] ),
    .A1(net3002),
    .S(net3173),
    .X(_01053_));
 sg13g2_mux2_1 _11042_ (.A0(\cpu.regs[6][13] ),
    .A1(net3019),
    .S(net3173),
    .X(_01054_));
 sg13g2_nor2_1 _11043_ (.A(\cpu.regs[6][14] ),
    .B(net3176),
    .Y(_04993_));
 sg13g2_a21oi_1 _11044_ (.A1(net3035),
    .A2(net3176),
    .Y(_01055_),
    .B1(_04993_));
 sg13g2_nor2_1 _11045_ (.A(\cpu.regs[6][15] ),
    .B(net3176),
    .Y(_04994_));
 sg13g2_a21oi_1 _11046_ (.A1(net3033),
    .A2(net3176),
    .Y(_01056_),
    .B1(_04994_));
 sg13g2_mux2_1 _11047_ (.A0(\cpu.regs[6][16] ),
    .A1(net2999),
    .S(net3173),
    .X(_01057_));
 sg13g2_nor2_1 _11048_ (.A(\cpu.regs[6][17] ),
    .B(net3177),
    .Y(_04995_));
 sg13g2_a21oi_1 _11049_ (.A1(net2997),
    .A2(net3177),
    .Y(_01058_),
    .B1(_04995_));
 sg13g2_mux2_1 _11050_ (.A0(\cpu.regs[6][18] ),
    .A1(net2995),
    .S(net3175),
    .X(_01059_));
 sg13g2_nor2_1 _11051_ (.A(\cpu.regs[6][19] ),
    .B(net3177),
    .Y(_04996_));
 sg13g2_a21oi_1 _11052_ (.A1(net2993),
    .A2(net3177),
    .Y(_01060_),
    .B1(_04996_));
 sg13g2_mux2_1 _11053_ (.A0(\cpu.regs[6][20] ),
    .A1(net2992),
    .S(net3173),
    .X(_01061_));
 sg13g2_mux2_1 _11054_ (.A0(\cpu.regs[6][21] ),
    .A1(net2990),
    .S(net3178),
    .X(_01062_));
 sg13g2_mux2_1 _11055_ (.A0(\cpu.regs[6][22] ),
    .A1(net3018),
    .S(net3175),
    .X(_01063_));
 sg13g2_mux2_1 _11056_ (.A0(\cpu.regs[6][23] ),
    .A1(net3015),
    .S(net3175),
    .X(_01064_));
 sg13g2_mux2_1 _11057_ (.A0(\cpu.regs[6][24] ),
    .A1(net2988),
    .S(net3175),
    .X(_01065_));
 sg13g2_mux2_1 _11058_ (.A0(\cpu.regs[6][25] ),
    .A1(net2985),
    .S(net3175),
    .X(_01066_));
 sg13g2_mux2_1 _11059_ (.A0(\cpu.regs[6][26] ),
    .A1(net3013),
    .S(net3173),
    .X(_01067_));
 sg13g2_mux2_1 _11060_ (.A0(\cpu.regs[6][27] ),
    .A1(net3011),
    .S(net3175),
    .X(_01068_));
 sg13g2_mux2_1 _11061_ (.A0(\cpu.regs[6][28] ),
    .A1(net2984),
    .S(net3175),
    .X(_01069_));
 sg13g2_mux2_1 _11062_ (.A0(\cpu.regs[6][29] ),
    .A1(net2981),
    .S(net3175),
    .X(_01070_));
 sg13g2_mux2_1 _11063_ (.A0(\cpu.regs[6][30] ),
    .A1(net3009),
    .S(net3173),
    .X(_01071_));
 sg13g2_mux2_1 _11064_ (.A0(\cpu.regs[6][31] ),
    .A1(net3007),
    .S(net3173),
    .X(_01072_));
 sg13g2_and2_2 _11065_ (.A(_04113_),
    .B(_04917_),
    .X(_04997_));
 sg13g2_mux2_1 _11066_ (.A0(\cpu.regs[5][0] ),
    .A1(net3046),
    .S(net3168),
    .X(_01073_));
 sg13g2_mux2_1 _11067_ (.A0(\cpu.regs[5][1] ),
    .A1(net3041),
    .S(net3168),
    .X(_01074_));
 sg13g2_mux2_1 _11068_ (.A0(\cpu.regs[5][2] ),
    .A1(net3040),
    .S(net3168),
    .X(_01075_));
 sg13g2_mux2_1 _11069_ (.A0(\cpu.regs[5][3] ),
    .A1(net3005),
    .S(net3170),
    .X(_01076_));
 sg13g2_mux2_1 _11070_ (.A0(\cpu.regs[5][4] ),
    .A1(net3003),
    .S(net3167),
    .X(_01077_));
 sg13g2_mux2_1 _11071_ (.A0(\cpu.regs[5][5] ),
    .A1(net3029),
    .S(net3171),
    .X(_01078_));
 sg13g2_mux2_1 _11072_ (.A0(\cpu.regs[5][6] ),
    .A1(net3037),
    .S(net3168),
    .X(_01079_));
 sg13g2_mux2_1 _11073_ (.A0(\cpu.regs[5][7] ),
    .A1(net3044),
    .S(net3170),
    .X(_01080_));
 sg13g2_mux2_1 _11074_ (.A0(\cpu.regs[5][8] ),
    .A1(net3027),
    .S(net3170),
    .X(_01081_));
 sg13g2_mux2_1 _11075_ (.A0(\cpu.regs[5][9] ),
    .A1(net3026),
    .S(net3170),
    .X(_01082_));
 sg13g2_mux2_1 _11076_ (.A0(\cpu.regs[5][10] ),
    .A1(net3023),
    .S(net3171),
    .X(_01083_));
 sg13g2_mux2_1 _11077_ (.A0(\cpu.regs[5][11] ),
    .A1(net3021),
    .S(net3171),
    .X(_01084_));
 sg13g2_mux2_1 _11078_ (.A0(\cpu.regs[5][12] ),
    .A1(net3002),
    .S(net3167),
    .X(_01085_));
 sg13g2_mux2_1 _11079_ (.A0(\cpu.regs[5][13] ),
    .A1(net3019),
    .S(net3167),
    .X(_01086_));
 sg13g2_nor2_1 _11080_ (.A(\cpu.regs[5][14] ),
    .B(net3170),
    .Y(_04998_));
 sg13g2_a21oi_1 _11081_ (.A1(net3035),
    .A2(net3170),
    .Y(_01087_),
    .B1(_04998_));
 sg13g2_nor2_1 _11082_ (.A(\cpu.regs[5][15] ),
    .B(net3170),
    .Y(_04999_));
 sg13g2_a21oi_1 _11083_ (.A1(net3033),
    .A2(net3170),
    .Y(_01088_),
    .B1(_04999_));
 sg13g2_mux2_1 _11084_ (.A0(\cpu.regs[5][16] ),
    .A1(net2999),
    .S(net3167),
    .X(_01089_));
 sg13g2_nor2_1 _11085_ (.A(\cpu.regs[5][17] ),
    .B(net3171),
    .Y(_05000_));
 sg13g2_a21oi_1 _11086_ (.A1(net2997),
    .A2(net3171),
    .Y(_01090_),
    .B1(_05000_));
 sg13g2_mux2_1 _11087_ (.A0(\cpu.regs[5][18] ),
    .A1(net2995),
    .S(net3169),
    .X(_01091_));
 sg13g2_nor2_1 _11088_ (.A(\cpu.regs[5][19] ),
    .B(net3169),
    .Y(_05001_));
 sg13g2_a21oi_1 _11089_ (.A1(net2993),
    .A2(net3169),
    .Y(_01092_),
    .B1(_05001_));
 sg13g2_mux2_1 _11090_ (.A0(\cpu.regs[5][20] ),
    .A1(net2992),
    .S(net3167),
    .X(_01093_));
 sg13g2_mux2_1 _11091_ (.A0(\cpu.regs[5][21] ),
    .A1(net2989),
    .S(net3172),
    .X(_01094_));
 sg13g2_mux2_1 _11092_ (.A0(\cpu.regs[5][22] ),
    .A1(net3018),
    .S(net3169),
    .X(_01095_));
 sg13g2_mux2_1 _11093_ (.A0(\cpu.regs[5][23] ),
    .A1(net3016),
    .S(net3172),
    .X(_01096_));
 sg13g2_mux2_1 _11094_ (.A0(\cpu.regs[5][24] ),
    .A1(net2988),
    .S(net3169),
    .X(_01097_));
 sg13g2_mux2_1 _11095_ (.A0(\cpu.regs[5][25] ),
    .A1(net2985),
    .S(net3172),
    .X(_01098_));
 sg13g2_mux2_1 _11096_ (.A0(\cpu.regs[5][26] ),
    .A1(net3013),
    .S(net3167),
    .X(_01099_));
 sg13g2_mux2_1 _11097_ (.A0(\cpu.regs[5][27] ),
    .A1(net3011),
    .S(net3169),
    .X(_01100_));
 sg13g2_mux2_1 _11098_ (.A0(\cpu.regs[5][28] ),
    .A1(net2984),
    .S(net3169),
    .X(_01101_));
 sg13g2_mux2_1 _11099_ (.A0(\cpu.regs[5][29] ),
    .A1(net2981),
    .S(net3169),
    .X(_01102_));
 sg13g2_mux2_1 _11100_ (.A0(\cpu.regs[5][30] ),
    .A1(net3009),
    .S(net3167),
    .X(_01103_));
 sg13g2_mux2_1 _11101_ (.A0(\cpu.regs[5][31] ),
    .A1(net3007),
    .S(net3167),
    .X(_01104_));
 sg13g2_nor3_2 _11102_ (.A(_02520_),
    .B(net3124),
    .C(_04867_),
    .Y(_05002_));
 sg13g2_mux2_1 _11103_ (.A0(\irqen[0] ),
    .A1(_02498_),
    .S(_05002_),
    .X(_01114_));
 sg13g2_mux2_1 _11104_ (.A0(\irqen[1] ),
    .A1(_02469_),
    .S(_05002_),
    .X(_01115_));
 sg13g2_mux2_1 _11105_ (.A0(\irqen[2] ),
    .A1(net3326),
    .S(_05002_),
    .X(_01116_));
 sg13g2_mux2_1 _11106_ (.A0(\irqen[3] ),
    .A1(net3327),
    .S(_05002_),
    .X(_01117_));
 sg13g2_nor2_1 _11107_ (.A(\irqen[4] ),
    .B(_05002_),
    .Y(_05003_));
 sg13g2_a21oi_1 _11108_ (.A1(_02928_),
    .A2(_05002_),
    .Y(_01118_),
    .B1(_05003_));
 sg13g2_nand2_2 _11109_ (.Y(_05004_),
    .A(net3720),
    .B(_03406_));
 sg13g2_mux2_1 _11110_ (.A0(\pwm[0] ),
    .A1(\pwmbuf[0] ),
    .S(_05004_),
    .X(_01119_));
 sg13g2_mux2_1 _11111_ (.A0(\pwm[1] ),
    .A1(\pwmbuf[1] ),
    .S(_05004_),
    .X(_01120_));
 sg13g2_mux2_1 _11112_ (.A0(\pwm[2] ),
    .A1(\pwmbuf[2] ),
    .S(_05004_),
    .X(_01121_));
 sg13g2_mux2_1 _11113_ (.A0(\pwm[3] ),
    .A1(\pwmbuf[3] ),
    .S(_05004_),
    .X(_01122_));
 sg13g2_mux2_1 _11114_ (.A0(\pwm[4] ),
    .A1(\pwmbuf[4] ),
    .S(_05004_),
    .X(_01123_));
 sg13g2_mux2_1 _11115_ (.A0(\pwm[5] ),
    .A1(\pwmbuf[5] ),
    .S(_05004_),
    .X(_01124_));
 sg13g2_mux2_1 _11116_ (.A0(\pwm[6] ),
    .A1(\pwmbuf[6] ),
    .S(_05004_),
    .X(_01125_));
 sg13g2_mux2_1 _11117_ (.A0(\pwm[7] ),
    .A1(\pwmbuf[7] ),
    .S(_05004_),
    .X(_01126_));
 sg13g2_nand3_1 _11118_ (.B(_02519_),
    .C(_03422_),
    .A(net3098),
    .Y(_05005_));
 sg13g2_nor2_1 _11119_ (.A(net3876),
    .B(_05005_),
    .Y(_05006_));
 sg13g2_mux2_1 _11120_ (.A0(\pwm[0] ),
    .A1(_02498_),
    .S(_05006_),
    .X(_01127_));
 sg13g2_mux2_1 _11121_ (.A0(\pwm[1] ),
    .A1(_02469_),
    .S(net3061),
    .X(_01128_));
 sg13g2_mux2_1 _11122_ (.A0(\pwm[2] ),
    .A1(_03101_),
    .S(net3061),
    .X(_01129_));
 sg13g2_mux2_1 _11123_ (.A0(\pwm[3] ),
    .A1(_03014_),
    .S(net3061),
    .X(_01130_));
 sg13g2_nor2_1 _11124_ (.A(\pwm[4] ),
    .B(net3061),
    .Y(_05007_));
 sg13g2_a21oi_1 _11125_ (.A1(_02928_),
    .A2(net3061),
    .Y(_01131_),
    .B1(_05007_));
 sg13g2_mux2_1 _11126_ (.A0(\pwm[5] ),
    .A1(_02842_),
    .S(net3061),
    .X(_01132_));
 sg13g2_mux2_1 _11127_ (.A0(\pwm[6] ),
    .A1(_02759_),
    .S(net3061),
    .X(_01133_));
 sg13g2_mux2_1 _11128_ (.A0(\pwm[7] ),
    .A1(net3330),
    .S(net3061),
    .X(_01134_));
 sg13g2_nor4_1 _11129_ (.A(\pwmc[5] ),
    .B(\pwmc[4] ),
    .C(\pwmc[7] ),
    .D(\pwmc[6] ),
    .Y(_05008_));
 sg13g2_nor4_1 _11130_ (.A(\pwmc[1] ),
    .B(\pwmc[0] ),
    .C(\pwmc[3] ),
    .D(\pwmc[2] ),
    .Y(_05009_));
 sg13g2_nand2_2 _11131_ (.Y(_05010_),
    .A(_05008_),
    .B(_05009_));
 sg13g2_nand2b_1 _11132_ (.Y(_05011_),
    .B(\pwmc[1] ),
    .A_N(\pwmbuf[1] ));
 sg13g2_xnor2_1 _11133_ (.Y(_05012_),
    .A(\pwmc[0] ),
    .B(\pwmbuf[0] ));
 sg13g2_xor2_1 _11134_ (.B(\pwmbuf[2] ),
    .A(\pwmc[2] ),
    .X(_05013_));
 sg13g2_nand2b_1 _11135_ (.Y(_05014_),
    .B(\pwmc[7] ),
    .A_N(\pwmbuf[7] ));
 sg13g2_nand2b_1 _11136_ (.Y(_05015_),
    .B(\pwmc[5] ),
    .A_N(\pwmbuf[5] ));
 sg13g2_nand2b_1 _11137_ (.Y(_05016_),
    .B(\pwmbuf[7] ),
    .A_N(\pwmc[7] ));
 sg13g2_xor2_1 _11138_ (.B(\pwmbuf[4] ),
    .A(\pwmc[4] ),
    .X(_05017_));
 sg13g2_a22oi_1 _11139_ (.Y(_05018_),
    .B1(\pwmbuf[5] ),
    .B2(_01704_),
    .A2(\pwmbuf[1] ),
    .A1(_01702_));
 sg13g2_xnor2_1 _11140_ (.Y(_05019_),
    .A(\pwmc[3] ),
    .B(\pwmbuf[3] ));
 sg13g2_xnor2_1 _11141_ (.Y(_05020_),
    .A(\pwmc[6] ),
    .B(\pwmbuf[6] ));
 sg13g2_nand4_1 _11142_ (.B(_05018_),
    .C(_05019_),
    .A(_05012_),
    .Y(_05021_),
    .D(_05020_));
 sg13g2_nand4_1 _11143_ (.B(_05014_),
    .C(_05015_),
    .A(_05011_),
    .Y(_05022_),
    .D(_05016_));
 sg13g2_nor4_1 _11144_ (.A(_05013_),
    .B(_05017_),
    .C(_05021_),
    .D(_05022_),
    .Y(_05023_));
 sg13g2_a21oi_1 _11145_ (.A1(_01706_),
    .A2(_05010_),
    .Y(_01135_),
    .B1(_05023_));
 sg13g2_nand3_1 _11146_ (.B(_02519_),
    .C(_03421_),
    .A(net3098),
    .Y(_05024_));
 sg13g2_a21o_1 _11147_ (.A2(_05024_),
    .A1(udirty),
    .B1(_02521_),
    .X(_01136_));
 sg13g2_nand2_1 _11148_ (.Y(_05025_),
    .A(pwmirq),
    .B(_05005_));
 sg13g2_nand2_1 _11149_ (.Y(_01137_),
    .A(_05010_),
    .B(_05025_));
 sg13g2_mux2_1 _11150_ (.A0(net900),
    .A1(_03329_),
    .S(net3724),
    .X(_01138_));
 sg13g2_nand2_1 _11151_ (.Y(_05026_),
    .A(net3724),
    .B(_03325_));
 sg13g2_o21ai_1 _11152_ (.B1(_05026_),
    .Y(_01139_),
    .A1(_01734_),
    .A2(net3724));
 sg13g2_mux2_1 _11153_ (.A0(net901),
    .A1(_03321_),
    .S(_02707_),
    .X(_01140_));
 sg13g2_mux2_1 _11154_ (.A0(net904),
    .A1(_03317_),
    .S(_02707_),
    .X(_01141_));
 sg13g2_mux2_1 _11155_ (.A0(net899),
    .A1(_03314_),
    .S(net3724),
    .X(_01142_));
 sg13g2_nor2_1 _11156_ (.A(net897),
    .B(net3724),
    .Y(_05027_));
 sg13g2_a21oi_1 _11157_ (.A1(net3724),
    .A2(_03309_),
    .Y(_01143_),
    .B1(_05027_));
 sg13g2_mux2_1 _11158_ (.A0(net903),
    .A1(_03302_),
    .S(net3724),
    .X(_01144_));
 sg13g2_mux2_1 _11159_ (.A0(net895),
    .A1(_03299_),
    .S(_02707_),
    .X(_01145_));
 sg13g2_mux2_1 _11160_ (.A0(_03329_),
    .A1(net922),
    .S(net3457),
    .X(_01146_));
 sg13g2_mux2_1 _11161_ (.A0(_03325_),
    .A1(net916),
    .S(_02705_),
    .X(_01147_));
 sg13g2_mux2_1 _11162_ (.A0(_03321_),
    .A1(net906),
    .S(net3457),
    .X(_01148_));
 sg13g2_mux2_1 _11163_ (.A0(_03317_),
    .A1(net909),
    .S(net3457),
    .X(_01149_));
 sg13g2_mux2_1 _11164_ (.A0(_03314_),
    .A1(net908),
    .S(_02705_),
    .X(_01150_));
 sg13g2_nand2_1 _11165_ (.Y(_05028_),
    .A(net891),
    .B(net3457));
 sg13g2_o21ai_1 _11166_ (.B1(_05028_),
    .Y(_01151_),
    .A1(net3457),
    .A2(_03309_));
 sg13g2_mux2_1 _11167_ (.A0(_03302_),
    .A1(net926),
    .S(net3457),
    .X(_01152_));
 sg13g2_mux2_1 _11168_ (.A0(_03299_),
    .A1(net919),
    .S(net3457),
    .X(_01153_));
 sg13g2_nand2_1 _11169_ (.Y(_05029_),
    .A(_04904_),
    .B(_04910_));
 sg13g2_mux2_1 _11170_ (.A0(net3047),
    .A1(\cpu.regs[8][0] ),
    .S(net3165),
    .X(_01154_));
 sg13g2_mux2_1 _11171_ (.A0(net3042),
    .A1(\cpu.regs[8][1] ),
    .S(net3165),
    .X(_01155_));
 sg13g2_mux2_1 _11172_ (.A0(net3039),
    .A1(\cpu.regs[8][2] ),
    .S(net3165),
    .X(_01156_));
 sg13g2_mux2_1 _11173_ (.A0(net3006),
    .A1(\cpu.regs[8][3] ),
    .S(net3164),
    .X(_01157_));
 sg13g2_mux2_1 _11174_ (.A0(net3004),
    .A1(\cpu.regs[8][4] ),
    .S(net3165),
    .X(_01158_));
 sg13g2_mux2_1 _11175_ (.A0(net3030),
    .A1(\cpu.regs[8][5] ),
    .S(net3164),
    .X(_01159_));
 sg13g2_mux2_1 _11176_ (.A0(net3037),
    .A1(\cpu.regs[8][6] ),
    .S(net3165),
    .X(_01160_));
 sg13g2_mux2_1 _11177_ (.A0(net3045),
    .A1(\cpu.regs[8][7] ),
    .S(net3164),
    .X(_01161_));
 sg13g2_mux2_1 _11178_ (.A0(net3028),
    .A1(\cpu.regs[8][8] ),
    .S(net3164),
    .X(_01162_));
 sg13g2_mux2_1 _11179_ (.A0(net3025),
    .A1(\cpu.regs[8][9] ),
    .S(net3165),
    .X(_01163_));
 sg13g2_mux2_1 _11180_ (.A0(net3024),
    .A1(\cpu.regs[8][10] ),
    .S(net3164),
    .X(_01164_));
 sg13g2_mux2_1 _11181_ (.A0(net3022),
    .A1(\cpu.regs[8][11] ),
    .S(net3163),
    .X(_01165_));
 sg13g2_mux2_1 _11182_ (.A0(net3002),
    .A1(\cpu.regs[8][12] ),
    .S(net3162),
    .X(_01166_));
 sg13g2_mux2_1 _11183_ (.A0(net3020),
    .A1(\cpu.regs[8][13] ),
    .S(net3162),
    .X(_01167_));
 sg13g2_nand2_1 _11184_ (.Y(_05030_),
    .A(\cpu.regs[8][14] ),
    .B(net3163));
 sg13g2_o21ai_1 _11185_ (.B1(_05030_),
    .Y(_01168_),
    .A1(net3036),
    .A2(net3163));
 sg13g2_nand2_1 _11186_ (.Y(_05031_),
    .A(\cpu.regs[8][15] ),
    .B(net3163));
 sg13g2_o21ai_1 _11187_ (.B1(_05031_),
    .Y(_01169_),
    .A1(net3034),
    .A2(net3163));
 sg13g2_mux2_1 _11188_ (.A0(net3000),
    .A1(\cpu.regs[8][16] ),
    .S(net3165),
    .X(_01170_));
 sg13g2_nand2_1 _11189_ (.Y(_05032_),
    .A(\cpu.regs[8][17] ),
    .B(net3163));
 sg13g2_o21ai_1 _11190_ (.B1(_05032_),
    .Y(_01171_),
    .A1(net2998),
    .A2(net3163));
 sg13g2_mux2_1 _11191_ (.A0(net2996),
    .A1(\cpu.regs[8][18] ),
    .S(net3163),
    .X(_01172_));
 sg13g2_nand2_1 _11192_ (.Y(_05033_),
    .A(\cpu.regs[8][19] ),
    .B(net3161));
 sg13g2_o21ai_1 _11193_ (.B1(_05033_),
    .Y(_01173_),
    .A1(net2994),
    .A2(net3161));
 sg13g2_mux2_1 _11194_ (.A0(net2991),
    .A1(\cpu.regs[8][20] ),
    .S(net3162),
    .X(_01174_));
 sg13g2_mux2_1 _11195_ (.A0(net2989),
    .A1(\cpu.regs[8][21] ),
    .S(net3161),
    .X(_01175_));
 sg13g2_mux2_1 _11196_ (.A0(net3017),
    .A1(\cpu.regs[8][22] ),
    .S(net3161),
    .X(_01176_));
 sg13g2_mux2_1 _11197_ (.A0(net3016),
    .A1(\cpu.regs[8][23] ),
    .S(net3161),
    .X(_01177_));
 sg13g2_mux2_1 _11198_ (.A0(net2987),
    .A1(\cpu.regs[8][24] ),
    .S(net3161),
    .X(_01178_));
 sg13g2_mux2_1 _11199_ (.A0(net2986),
    .A1(\cpu.regs[8][25] ),
    .S(net3161),
    .X(_01179_));
 sg13g2_mux2_1 _11200_ (.A0(net3014),
    .A1(\cpu.regs[8][26] ),
    .S(net3162),
    .X(_01180_));
 sg13g2_mux2_1 _11201_ (.A0(net3012),
    .A1(\cpu.regs[8][27] ),
    .S(net3161),
    .X(_01181_));
 sg13g2_mux2_1 _11202_ (.A0(net2983),
    .A1(\cpu.regs[8][28] ),
    .S(net3162),
    .X(_01182_));
 sg13g2_mux2_1 _11203_ (.A0(net2982),
    .A1(\cpu.regs[8][29] ),
    .S(net3166),
    .X(_01183_));
 sg13g2_mux2_1 _11204_ (.A0(net3010),
    .A1(\cpu.regs[8][30] ),
    .S(net3162),
    .X(_01184_));
 sg13g2_mux2_1 _11205_ (.A0(net3008),
    .A1(\cpu.regs[8][31] ),
    .S(net3162),
    .X(_01185_));
 sg13g2_nand4_1 _11206_ (.B(\cpu.Bimm[11] ),
    .C(net3701),
    .A(\cpu.Bimm[1] ),
    .Y(_05034_),
    .D(_04124_));
 sg13g2_mux2_1 _11207_ (.A0(net3047),
    .A1(\cpu.regs[15][0] ),
    .S(net3160),
    .X(_01186_));
 sg13g2_mux2_1 _11208_ (.A0(net3042),
    .A1(\cpu.regs[15][1] ),
    .S(net3160),
    .X(_01187_));
 sg13g2_mux2_1 _11209_ (.A0(net3039),
    .A1(\cpu.regs[15][2] ),
    .S(net3160),
    .X(_01188_));
 sg13g2_mux2_1 _11210_ (.A0(net3006),
    .A1(\cpu.regs[15][3] ),
    .S(net3159),
    .X(_01189_));
 sg13g2_mux2_1 _11211_ (.A0(net3004),
    .A1(\cpu.regs[15][4] ),
    .S(net3160),
    .X(_01190_));
 sg13g2_mux2_1 _11212_ (.A0(net3030),
    .A1(\cpu.regs[15][5] ),
    .S(net3159),
    .X(_01191_));
 sg13g2_mux2_1 _11213_ (.A0(net3038),
    .A1(\cpu.regs[15][6] ),
    .S(net3160),
    .X(_01192_));
 sg13g2_mux2_1 _11214_ (.A0(net3045),
    .A1(\cpu.regs[15][7] ),
    .S(net3159),
    .X(_01193_));
 sg13g2_mux2_1 _11215_ (.A0(net3027),
    .A1(\cpu.regs[15][8] ),
    .S(net3158),
    .X(_01194_));
 sg13g2_mux2_1 _11216_ (.A0(net3025),
    .A1(\cpu.regs[15][9] ),
    .S(net3159),
    .X(_01195_));
 sg13g2_mux2_1 _11217_ (.A0(net3024),
    .A1(\cpu.regs[15][10] ),
    .S(net3158),
    .X(_01196_));
 sg13g2_mux2_1 _11218_ (.A0(net3022),
    .A1(\cpu.regs[15][11] ),
    .S(net3158),
    .X(_01197_));
 sg13g2_mux2_1 _11219_ (.A0(net3001),
    .A1(\cpu.regs[15][12] ),
    .S(net3157),
    .X(_01198_));
 sg13g2_mux2_1 _11220_ (.A0(net3020),
    .A1(\cpu.regs[15][13] ),
    .S(net3157),
    .X(_01199_));
 sg13g2_nand2_1 _11221_ (.Y(_05035_),
    .A(\cpu.regs[15][14] ),
    .B(net3159));
 sg13g2_o21ai_1 _11222_ (.B1(_05035_),
    .Y(_01200_),
    .A1(net3036),
    .A2(net3159));
 sg13g2_nand2_1 _11223_ (.Y(_05036_),
    .A(\cpu.regs[15][15] ),
    .B(net3158));
 sg13g2_o21ai_1 _11224_ (.B1(_05036_),
    .Y(_01201_),
    .A1(net3034),
    .A2(net3158));
 sg13g2_mux2_1 _11225_ (.A0(net3000),
    .A1(\cpu.regs[15][16] ),
    .S(net3160),
    .X(_01202_));
 sg13g2_nand2_1 _11226_ (.Y(_05037_),
    .A(\cpu.regs[15][17] ),
    .B(net3158));
 sg13g2_o21ai_1 _11227_ (.B1(_05037_),
    .Y(_01203_),
    .A1(net2998),
    .A2(net3158));
 sg13g2_mux2_1 _11228_ (.A0(net2996),
    .A1(\cpu.regs[15][18] ),
    .S(net3155),
    .X(_01204_));
 sg13g2_nand2_1 _11229_ (.Y(_05038_),
    .A(\cpu.regs[15][19] ),
    .B(net3156));
 sg13g2_o21ai_1 _11230_ (.B1(_05038_),
    .Y(_01205_),
    .A1(net2994),
    .A2(net3156));
 sg13g2_mux2_1 _11231_ (.A0(net2991),
    .A1(\cpu.regs[15][20] ),
    .S(net3157),
    .X(_01206_));
 sg13g2_mux2_1 _11232_ (.A0(net2990),
    .A1(\cpu.regs[15][21] ),
    .S(net3155),
    .X(_01207_));
 sg13g2_mux2_1 _11233_ (.A0(net3017),
    .A1(\cpu.regs[15][22] ),
    .S(net3155),
    .X(_01208_));
 sg13g2_mux2_1 _11234_ (.A0(net3015),
    .A1(\cpu.regs[15][23] ),
    .S(net3155),
    .X(_01209_));
 sg13g2_mux2_1 _11235_ (.A0(net2988),
    .A1(\cpu.regs[15][24] ),
    .S(net3155),
    .X(_01210_));
 sg13g2_mux2_1 _11236_ (.A0(net2985),
    .A1(\cpu.regs[15][25] ),
    .S(net3155),
    .X(_01211_));
 sg13g2_mux2_1 _11237_ (.A0(net3014),
    .A1(\cpu.regs[15][26] ),
    .S(net3155),
    .X(_01212_));
 sg13g2_mux2_1 _11238_ (.A0(net3012),
    .A1(\cpu.regs[15][27] ),
    .S(net3156),
    .X(_01213_));
 sg13g2_mux2_1 _11239_ (.A0(net2983),
    .A1(\cpu.regs[15][28] ),
    .S(net3156),
    .X(_01214_));
 sg13g2_mux2_1 _11240_ (.A0(net2981),
    .A1(\cpu.regs[15][29] ),
    .S(net3158),
    .X(_01215_));
 sg13g2_mux2_1 _11241_ (.A0(net3010),
    .A1(\cpu.regs[15][30] ),
    .S(net3157),
    .X(_01216_));
 sg13g2_mux2_1 _11242_ (.A0(net3008),
    .A1(\cpu.regs[15][31] ),
    .S(net3155),
    .X(_01217_));
 sg13g2_and2_1 _11243_ (.A(_04113_),
    .B(_04904_),
    .X(_05039_));
 sg13g2_mux2_1 _11244_ (.A0(\cpu.regs[9][0] ),
    .A1(net3046),
    .S(net3153),
    .X(_01218_));
 sg13g2_mux2_1 _11245_ (.A0(\cpu.regs[9][1] ),
    .A1(net3042),
    .S(net3153),
    .X(_01219_));
 sg13g2_mux2_1 _11246_ (.A0(\cpu.regs[9][2] ),
    .A1(net3039),
    .S(net3153),
    .X(_01220_));
 sg13g2_mux2_1 _11247_ (.A0(\cpu.regs[9][3] ),
    .A1(net3005),
    .S(net3152),
    .X(_01221_));
 sg13g2_mux2_1 _11248_ (.A0(\cpu.regs[9][4] ),
    .A1(net3004),
    .S(net3153),
    .X(_01222_));
 sg13g2_mux2_1 _11249_ (.A0(\cpu.regs[9][5] ),
    .A1(net3029),
    .S(net3152),
    .X(_01223_));
 sg13g2_mux2_1 _11250_ (.A0(\cpu.regs[9][6] ),
    .A1(net3037),
    .S(net3153),
    .X(_01224_));
 sg13g2_mux2_1 _11251_ (.A0(\cpu.regs[9][7] ),
    .A1(net3044),
    .S(net3152),
    .X(_01225_));
 sg13g2_mux2_1 _11252_ (.A0(\cpu.regs[9][8] ),
    .A1(net3028),
    .S(net3151),
    .X(_01226_));
 sg13g2_mux2_1 _11253_ (.A0(\cpu.regs[9][9] ),
    .A1(net3025),
    .S(net3153),
    .X(_01227_));
 sg13g2_mux2_1 _11254_ (.A0(\cpu.regs[9][10] ),
    .A1(net3023),
    .S(net3152),
    .X(_01228_));
 sg13g2_mux2_1 _11255_ (.A0(\cpu.regs[9][11] ),
    .A1(net3021),
    .S(net3151),
    .X(_01229_));
 sg13g2_mux2_1 _11256_ (.A0(\cpu.regs[9][12] ),
    .A1(net3001),
    .S(net3150),
    .X(_01230_));
 sg13g2_mux2_1 _11257_ (.A0(\cpu.regs[9][13] ),
    .A1(net3019),
    .S(net3150),
    .X(_01231_));
 sg13g2_nor2_1 _11258_ (.A(\cpu.regs[9][14] ),
    .B(net3151),
    .Y(_05040_));
 sg13g2_a21oi_1 _11259_ (.A1(net3035),
    .A2(net3151),
    .Y(_01232_),
    .B1(_05040_));
 sg13g2_nor2_1 _11260_ (.A(\cpu.regs[9][15] ),
    .B(net3151),
    .Y(_05041_));
 sg13g2_a21oi_1 _11261_ (.A1(net3033),
    .A2(net3151),
    .Y(_01233_),
    .B1(_05041_));
 sg13g2_mux2_1 _11262_ (.A0(\cpu.regs[9][16] ),
    .A1(net2999),
    .S(net3153),
    .X(_01234_));
 sg13g2_nor2_1 _11263_ (.A(\cpu.regs[9][17] ),
    .B(net3151),
    .Y(_05042_));
 sg13g2_a21oi_1 _11264_ (.A1(net2997),
    .A2(net3151),
    .Y(_01235_),
    .B1(_05042_));
 sg13g2_mux2_1 _11265_ (.A0(\cpu.regs[9][18] ),
    .A1(net2995),
    .S(net3154),
    .X(_01236_));
 sg13g2_nor2_1 _11266_ (.A(\cpu.regs[9][19] ),
    .B(net3149),
    .Y(_05043_));
 sg13g2_a21oi_1 _11267_ (.A1(net2993),
    .A2(net3149),
    .Y(_01237_),
    .B1(_05043_));
 sg13g2_mux2_1 _11268_ (.A0(\cpu.regs[9][20] ),
    .A1(net2991),
    .S(net3150),
    .X(_01238_));
 sg13g2_mux2_1 _11269_ (.A0(\cpu.regs[9][21] ),
    .A1(net2989),
    .S(net3149),
    .X(_01239_));
 sg13g2_mux2_1 _11270_ (.A0(\cpu.regs[9][22] ),
    .A1(net3017),
    .S(net3149),
    .X(_01240_));
 sg13g2_mux2_1 _11271_ (.A0(\cpu.regs[9][23] ),
    .A1(net3016),
    .S(net3149),
    .X(_01241_));
 sg13g2_mux2_1 _11272_ (.A0(\cpu.regs[9][24] ),
    .A1(net2987),
    .S(net3149),
    .X(_01242_));
 sg13g2_mux2_1 _11273_ (.A0(\cpu.regs[9][25] ),
    .A1(net2986),
    .S(net3154),
    .X(_01243_));
 sg13g2_mux2_1 _11274_ (.A0(\cpu.regs[9][26] ),
    .A1(net3014),
    .S(net3150),
    .X(_01244_));
 sg13g2_mux2_1 _11275_ (.A0(\cpu.regs[9][27] ),
    .A1(net3012),
    .S(net3149),
    .X(_01245_));
 sg13g2_mux2_1 _11276_ (.A0(\cpu.regs[9][28] ),
    .A1(net2983),
    .S(net3150),
    .X(_01246_));
 sg13g2_mux2_1 _11277_ (.A0(\cpu.regs[9][29] ),
    .A1(net2982),
    .S(net3149),
    .X(_01247_));
 sg13g2_mux2_1 _11278_ (.A0(\cpu.regs[9][30] ),
    .A1(net3010),
    .S(net3150),
    .X(_01248_));
 sg13g2_mux2_1 _11279_ (.A0(\cpu.regs[9][31] ),
    .A1(net3007),
    .S(net3150),
    .X(_01249_));
 sg13g2_nand2_1 _11280_ (.Y(_05044_),
    .A(\cpu.PCreg1[2] ),
    .B(_03355_));
 sg13g2_nor2_1 _11281_ (.A(net3627),
    .B(_04075_),
    .Y(_05045_));
 sg13g2_nand2_1 _11282_ (.Y(_05046_),
    .A(net3635),
    .B(_04074_));
 sg13g2_nand2_1 _11283_ (.Y(_05047_),
    .A(\cpu.IR[22] ),
    .B(net3415));
 sg13g2_o21ai_1 _11284_ (.B1(_05047_),
    .Y(_05048_),
    .A1(_00549_),
    .A2(net3115));
 sg13g2_nand2_1 _11285_ (.Y(_05049_),
    .A(_01725_),
    .B(_05048_));
 sg13g2_o21ai_1 _11286_ (.B1(net3108),
    .Y(_05050_),
    .A1(_01725_),
    .A2(_05048_));
 sg13g2_nand2b_1 _11287_ (.Y(_05051_),
    .B(_05049_),
    .A_N(_05050_));
 sg13g2_nor2b_1 _11288_ (.A(_04073_),
    .B_N(\cpu.PC[2] ),
    .Y(_05052_));
 sg13g2_xnor2_1 _11289_ (.Y(_05053_),
    .A(\cpu.PC[2] ),
    .B(_04073_));
 sg13g2_a21oi_1 _11290_ (.A1(net3113),
    .A2(_05053_),
    .Y(_05054_),
    .B1(net3424));
 sg13g2_a22oi_1 _11291_ (.Y(_05055_),
    .B1(_05051_),
    .B2(_05054_),
    .A2(_04024_),
    .A1(net3424));
 sg13g2_inv_1 _11292_ (.Y(_05056_),
    .A(_05055_));
 sg13g2_nor2_1 _11293_ (.A(net3309),
    .B(_05055_),
    .Y(_05057_));
 sg13g2_nor2b_1 _11294_ (.A(_04079_),
    .B_N(_04076_),
    .Y(_05058_));
 sg13g2_nor2_1 _11295_ (.A(_04071_),
    .B(_05058_),
    .Y(_05059_));
 sg13g2_mux4_1 _11296_ (.S0(net3323),
    .A0(\irqvect[0][0] ),
    .A1(\irqvect[2][0] ),
    .A2(\irqvect[1][0] ),
    .A3(\irqvect[3][0] ),
    .S1(net3248),
    .X(_05060_));
 sg13g2_o21ai_1 _11297_ (.B1(net3715),
    .Y(_05061_),
    .A1(net3259),
    .A2(_05060_));
 sg13g2_o21ai_1 _11298_ (.B1(_05044_),
    .Y(_01346_),
    .A1(_05057_),
    .A2(_05061_));
 sg13g2_xor2_1 _11299_ (.B(_05052_),
    .A(\cpu.PC[3] ),
    .X(_05062_));
 sg13g2_a21oi_1 _11300_ (.A1(net3113),
    .A2(_05062_),
    .Y(_05063_),
    .B1(net3423));
 sg13g2_nand2_1 _11301_ (.Y(_05064_),
    .A(\cpu.IR[23] ),
    .B(net3414));
 sg13g2_o21ai_1 _11302_ (.B1(_05064_),
    .Y(_05065_),
    .A1(_00550_),
    .A2(net3115));
 sg13g2_nand2_1 _11303_ (.Y(_05066_),
    .A(_01726_),
    .B(_05065_));
 sg13g2_xnor2_1 _11304_ (.Y(_05067_),
    .A(_01726_),
    .B(_05065_));
 sg13g2_xnor2_1 _11305_ (.Y(_05068_),
    .A(_05049_),
    .B(_05067_));
 sg13g2_o21ai_1 _11306_ (.B1(_05063_),
    .Y(_05069_),
    .A1(net3113),
    .A2(_05068_));
 sg13g2_o21ai_1 _11307_ (.B1(_05069_),
    .Y(_05070_),
    .A1(net3389),
    .A2(_04023_));
 sg13g2_mux4_1 _11308_ (.S0(net3323),
    .A0(\irqvect[0][1] ),
    .A1(\irqvect[2][1] ),
    .A2(\irqvect[1][1] ),
    .A3(\irqvect[3][1] ),
    .S1(net3249),
    .X(_05071_));
 sg13g2_o21ai_1 _11309_ (.B1(net3715),
    .Y(_05072_),
    .A1(net3258),
    .A2(_05071_));
 sg13g2_a21oi_1 _11310_ (.A1(net3259),
    .A2(_05070_),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_a21o_1 _11311_ (.A2(_03355_),
    .A1(\cpu.PCreg1[3] ),
    .B1(_05073_),
    .X(_01347_));
 sg13g2_nand2_1 _11312_ (.Y(_05074_),
    .A(\cpu.PCreg1[4] ),
    .B(net3876));
 sg13g2_o21ai_1 _11313_ (.B1(_05066_),
    .Y(_05075_),
    .A1(_05049_),
    .A2(_05067_));
 sg13g2_nand2_1 _11314_ (.Y(_05076_),
    .A(\cpu.IR[24] ),
    .B(net3414));
 sg13g2_o21ai_1 _11315_ (.B1(_05076_),
    .Y(_05077_),
    .A1(_00551_),
    .A2(net3115));
 sg13g2_xor2_1 _11316_ (.B(_05077_),
    .A(\cpu.PCci[4] ),
    .X(_05078_));
 sg13g2_nand2_1 _11317_ (.Y(_05079_),
    .A(_05075_),
    .B(_05078_));
 sg13g2_xor2_1 _11318_ (.B(_05078_),
    .A(_05075_),
    .X(_05080_));
 sg13g2_nand3_1 _11319_ (.B(\cpu.PC[3] ),
    .C(_05052_),
    .A(\cpu.PC[4] ),
    .Y(_05081_));
 sg13g2_a21o_1 _11320_ (.A2(_05052_),
    .A1(\cpu.PC[3] ),
    .B1(\cpu.PC[4] ),
    .X(_05082_));
 sg13g2_nand2_1 _11321_ (.Y(_05083_),
    .A(_05081_),
    .B(_05082_));
 sg13g2_o21ai_1 _11322_ (.B1(net3389),
    .Y(_05084_),
    .A1(net3108),
    .A2(_05083_));
 sg13g2_a21oi_1 _11323_ (.A1(net3107),
    .A2(_05080_),
    .Y(_05085_),
    .B1(_05084_));
 sg13g2_a21oi_2 _11324_ (.B1(_05085_),
    .Y(_05086_),
    .A2(_04027_),
    .A1(net3423));
 sg13g2_inv_1 _11325_ (.Y(_05087_),
    .A(_05086_));
 sg13g2_nor2_1 _11326_ (.A(net3309),
    .B(_05086_),
    .Y(_05088_));
 sg13g2_mux4_1 _11327_ (.S0(net3323),
    .A0(\irqvect[0][2] ),
    .A1(\irqvect[2][2] ),
    .A2(\irqvect[1][2] ),
    .A3(\irqvect[3][2] ),
    .S1(net3250),
    .X(_05089_));
 sg13g2_o21ai_1 _11328_ (.B1(net3706),
    .Y(_05090_),
    .A1(net3254),
    .A2(_05089_));
 sg13g2_o21ai_1 _11329_ (.B1(_05074_),
    .Y(_01348_),
    .A1(_05088_),
    .A2(_05090_));
 sg13g2_nand2_1 _11330_ (.Y(_05091_),
    .A(\cpu.Bimm[5] ),
    .B(net3414));
 sg13g2_o21ai_1 _11331_ (.B1(_05091_),
    .Y(_05092_),
    .A1(_00557_),
    .A2(net3115));
 sg13g2_nor2_1 _11332_ (.A(\cpu.PCci[5] ),
    .B(_05092_),
    .Y(_05093_));
 sg13g2_nand2_1 _11333_ (.Y(_05094_),
    .A(\cpu.PCci[5] ),
    .B(_05092_));
 sg13g2_xor2_1 _11334_ (.B(_05092_),
    .A(\cpu.PCci[5] ),
    .X(_05095_));
 sg13g2_nand2b_1 _11335_ (.Y(_05096_),
    .B(_05077_),
    .A_N(_00565_));
 sg13g2_nand2_1 _11336_ (.Y(_05097_),
    .A(_05079_),
    .B(_05096_));
 sg13g2_a21oi_1 _11337_ (.A1(_05095_),
    .A2(_05097_),
    .Y(_05098_),
    .B1(net3112));
 sg13g2_o21ai_1 _11338_ (.B1(_05098_),
    .Y(_05099_),
    .A1(_05095_),
    .A2(_05097_));
 sg13g2_nand2b_1 _11339_ (.Y(_05100_),
    .B(\cpu.PC[5] ),
    .A_N(_05081_));
 sg13g2_nand2b_1 _11340_ (.Y(_05101_),
    .B(_05081_),
    .A_N(\cpu.PC[5] ));
 sg13g2_nand3_1 _11341_ (.B(_05100_),
    .C(_05101_),
    .A(net3112),
    .Y(_05102_));
 sg13g2_a21oi_1 _11342_ (.A1(_05099_),
    .A2(_05102_),
    .Y(_05103_),
    .B1(net3423));
 sg13g2_a21oi_2 _11343_ (.B1(_05103_),
    .Y(_05104_),
    .A2(_04021_),
    .A1(net3423));
 sg13g2_mux4_1 _11344_ (.S0(net3323),
    .A0(\irqvect[0][3] ),
    .A1(\irqvect[2][3] ),
    .A2(\irqvect[1][3] ),
    .A3(\irqvect[3][3] ),
    .S1(net3249),
    .X(_05105_));
 sg13g2_o21ai_1 _11345_ (.B1(net3715),
    .Y(_05106_),
    .A1(net3258),
    .A2(_05105_));
 sg13g2_a21oi_1 _11346_ (.A1(net3259),
    .A2(_05104_),
    .Y(_05107_),
    .B1(_05106_));
 sg13g2_a21o_1 _11347_ (.A2(net3876),
    .A1(\cpu.PCreg1[5] ),
    .B1(_05107_),
    .X(_01349_));
 sg13g2_and2_1 _11348_ (.A(_05078_),
    .B(_05095_),
    .X(_05108_));
 sg13g2_o21ai_1 _11349_ (.B1(_05094_),
    .Y(_05109_),
    .A1(_05093_),
    .A2(_05096_));
 sg13g2_a21o_2 _11350_ (.A2(_05108_),
    .A1(_05075_),
    .B1(_05109_),
    .X(_05110_));
 sg13g2_nand2_1 _11351_ (.Y(_05111_),
    .A(\cpu.Bimm[6] ),
    .B(net3414));
 sg13g2_o21ai_1 _11352_ (.B1(_05111_),
    .Y(_05112_),
    .A1(_00558_),
    .A2(net3115));
 sg13g2_xor2_1 _11353_ (.B(_05112_),
    .A(\cpu.PCci[6] ),
    .X(_05113_));
 sg13g2_nand2_1 _11354_ (.Y(_05114_),
    .A(_05110_),
    .B(_05113_));
 sg13g2_xnor2_1 _11355_ (.Y(_05115_),
    .A(_05110_),
    .B(_05113_));
 sg13g2_nand2b_2 _11356_ (.Y(_05116_),
    .B(\cpu.PC[6] ),
    .A_N(_05100_));
 sg13g2_xnor2_1 _11357_ (.Y(_05117_),
    .A(\cpu.PC[6] ),
    .B(_05100_));
 sg13g2_a21oi_1 _11358_ (.A1(net3112),
    .A2(_05117_),
    .Y(_05118_),
    .B1(net3423));
 sg13g2_o21ai_1 _11359_ (.B1(_05118_),
    .Y(_05119_),
    .A1(net3112),
    .A2(_05115_));
 sg13g2_o21ai_1 _11360_ (.B1(_05119_),
    .Y(_05120_),
    .A1(net3389),
    .A2(_04018_));
 sg13g2_mux4_1 _11361_ (.S0(net3324),
    .A0(\irqvect[0][4] ),
    .A1(\irqvect[2][4] ),
    .A2(\irqvect[1][4] ),
    .A3(\irqvect[3][4] ),
    .S1(net3249),
    .X(_05121_));
 sg13g2_o21ai_1 _11362_ (.B1(net3714),
    .Y(_05122_),
    .A1(net3258),
    .A2(_05121_));
 sg13g2_a21oi_1 _11363_ (.A1(net3259),
    .A2(_05120_),
    .Y(_05123_),
    .B1(_05122_));
 sg13g2_a21o_1 _11364_ (.A2(net3876),
    .A1(\cpu.PCreg1[6] ),
    .B1(_05123_),
    .X(_01350_));
 sg13g2_nand2_1 _11365_ (.Y(_05124_),
    .A(\cpu.Bimm[7] ),
    .B(net3414));
 sg13g2_o21ai_1 _11366_ (.B1(_05124_),
    .Y(_05125_),
    .A1(_00559_),
    .A2(net3115));
 sg13g2_nor2_1 _11367_ (.A(\cpu.PCci[7] ),
    .B(_05125_),
    .Y(_05126_));
 sg13g2_nand2_1 _11368_ (.Y(_05127_),
    .A(\cpu.PCci[7] ),
    .B(_05125_));
 sg13g2_xor2_1 _11369_ (.B(_05125_),
    .A(\cpu.PCci[7] ),
    .X(_05128_));
 sg13g2_nand2b_1 _11370_ (.Y(_05129_),
    .B(_05112_),
    .A_N(_00566_));
 sg13g2_nand2_1 _11371_ (.Y(_05130_),
    .A(_05114_),
    .B(_05129_));
 sg13g2_o21ai_1 _11372_ (.B1(net3107),
    .Y(_05131_),
    .A1(_05128_),
    .A2(_05130_));
 sg13g2_a21oi_1 _11373_ (.A1(_05128_),
    .A2(_05130_),
    .Y(_05132_),
    .B1(_05131_));
 sg13g2_nand2b_1 _11374_ (.Y(_05133_),
    .B(\cpu.PC[7] ),
    .A_N(_05116_));
 sg13g2_xor2_1 _11375_ (.B(_05116_),
    .A(\cpu.PC[7] ),
    .X(_05134_));
 sg13g2_o21ai_1 _11376_ (.B1(net3389),
    .Y(_05135_),
    .A1(net3107),
    .A2(_05134_));
 sg13g2_nand2_1 _11377_ (.Y(_05136_),
    .A(net3424),
    .B(_04037_));
 sg13g2_o21ai_1 _11378_ (.B1(_05136_),
    .Y(_05137_),
    .A1(_05132_),
    .A2(_05135_));
 sg13g2_mux2_1 _11379_ (.A0(\irqvect[2][5] ),
    .A1(\irqvect[3][5] ),
    .S(net3250),
    .X(_05138_));
 sg13g2_mux2_1 _11380_ (.A0(\irqvect[0][5] ),
    .A1(\irqvect[1][5] ),
    .S(net3249),
    .X(_05139_));
 sg13g2_nand2_1 _11381_ (.Y(_05140_),
    .A(net3320),
    .B(_05139_));
 sg13g2_a21oi_1 _11382_ (.A1(net3323),
    .A2(_05138_),
    .Y(_05141_),
    .B1(net3258));
 sg13g2_a221oi_1 _11383_ (.B2(_05141_),
    .C1(net3875),
    .B1(_05140_),
    .A1(net3258),
    .Y(_05142_),
    .A2(_05137_));
 sg13g2_a21o_1 _11384_ (.A2(net3875),
    .A1(\cpu.PCreg1[7] ),
    .B1(_05142_),
    .X(_01351_));
 sg13g2_nand2b_1 _11385_ (.Y(_05143_),
    .B(\cpu.PC[8] ),
    .A_N(_05133_));
 sg13g2_xnor2_1 _11386_ (.Y(_05144_),
    .A(\cpu.PC[8] ),
    .B(_05133_));
 sg13g2_a21oi_1 _11387_ (.A1(net3112),
    .A2(_05144_),
    .Y(_05145_),
    .B1(net3424));
 sg13g2_o21ai_1 _11388_ (.B1(_05127_),
    .Y(_05146_),
    .A1(_05126_),
    .A2(_05129_));
 sg13g2_and2_1 _11389_ (.A(_05113_),
    .B(_05128_),
    .X(_05147_));
 sg13g2_a21oi_1 _11390_ (.A1(_05110_),
    .A2(_05147_),
    .Y(_05148_),
    .B1(_05146_));
 sg13g2_nand2_1 _11391_ (.Y(_05149_),
    .A(\cpu.Bimm[8] ),
    .B(net3414));
 sg13g2_o21ai_1 _11392_ (.B1(_05149_),
    .Y(_05150_),
    .A1(_00560_),
    .A2(net3115));
 sg13g2_xor2_1 _11393_ (.B(_05150_),
    .A(\cpu.PCci[8] ),
    .X(_05151_));
 sg13g2_nand2b_1 _11394_ (.Y(_05152_),
    .B(_05148_),
    .A_N(_05151_));
 sg13g2_nor2b_1 _11395_ (.A(_05148_),
    .B_N(_05151_),
    .Y(_05153_));
 sg13g2_nand2_1 _11396_ (.Y(_05154_),
    .A(net3107),
    .B(_05152_));
 sg13g2_o21ai_1 _11397_ (.B1(_05145_),
    .Y(_05155_),
    .A1(_05153_),
    .A2(_05154_));
 sg13g2_o21ai_1 _11398_ (.B1(_05155_),
    .Y(_05156_),
    .A1(net3389),
    .A2(_04019_));
 sg13g2_mux4_1 _11399_ (.S0(net3323),
    .A0(\irqvect[0][6] ),
    .A1(\irqvect[2][6] ),
    .A2(\irqvect[1][6] ),
    .A3(\irqvect[3][6] ),
    .S1(net3249),
    .X(_05157_));
 sg13g2_o21ai_1 _11400_ (.B1(net3706),
    .Y(_05158_),
    .A1(net3258),
    .A2(_05157_));
 sg13g2_a21oi_1 _11401_ (.A1(net3259),
    .A2(_05156_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_a21o_1 _11402_ (.A2(net3876),
    .A1(\cpu.PCreg1[8] ),
    .B1(_05159_),
    .X(_01352_));
 sg13g2_nand2_1 _11403_ (.Y(_05160_),
    .A(\cpu.PCreg1[9] ),
    .B(net3874));
 sg13g2_nand2_1 _11404_ (.Y(_05161_),
    .A(\cpu.Bimm[9] ),
    .B(net3414));
 sg13g2_o21ai_1 _11405_ (.B1(_05161_),
    .Y(_05162_),
    .A1(_00561_),
    .A2(net3115));
 sg13g2_nand2_1 _11406_ (.Y(_05163_),
    .A(\cpu.PCci[9] ),
    .B(_05162_));
 sg13g2_xor2_1 _11407_ (.B(_05162_),
    .A(\cpu.PCci[9] ),
    .X(_05164_));
 sg13g2_nor2b_1 _11408_ (.A(_00567_),
    .B_N(_05150_),
    .Y(_05165_));
 sg13g2_o21ai_1 _11409_ (.B1(_05164_),
    .Y(_05166_),
    .A1(_05153_),
    .A2(_05165_));
 sg13g2_or3_1 _11410_ (.A(_05153_),
    .B(_05164_),
    .C(_05165_),
    .X(_05167_));
 sg13g2_nand3_1 _11411_ (.B(_05166_),
    .C(_05167_),
    .A(net3107),
    .Y(_05168_));
 sg13g2_nor2b_1 _11412_ (.A(_05143_),
    .B_N(\cpu.PC[9] ),
    .Y(_05169_));
 sg13g2_xnor2_1 _11413_ (.Y(_05170_),
    .A(\cpu.PC[9] ),
    .B(_05143_));
 sg13g2_a21oi_1 _11414_ (.A1(net3112),
    .A2(_05170_),
    .Y(_05171_),
    .B1(net3424));
 sg13g2_a22oi_1 _11415_ (.Y(_05172_),
    .B1(_05168_),
    .B2(_05171_),
    .A2(_04030_),
    .A1(net3424));
 sg13g2_mux2_1 _11416_ (.A0(\irqvect[0][7] ),
    .A1(\irqvect[1][7] ),
    .S(net3249),
    .X(_05173_));
 sg13g2_nand2b_1 _11417_ (.Y(_05174_),
    .B(net3249),
    .A_N(\irqvect[3][7] ));
 sg13g2_o21ai_1 _11418_ (.B1(_05174_),
    .Y(_05175_),
    .A1(\irqvect[2][7] ),
    .A2(net3249));
 sg13g2_a21oi_1 _11419_ (.A1(net3319),
    .A2(_05173_),
    .Y(_05176_),
    .B1(net3258));
 sg13g2_o21ai_1 _11420_ (.B1(_05176_),
    .Y(_05177_),
    .A1(net3320),
    .A2(_05175_));
 sg13g2_o21ai_1 _11421_ (.B1(_05177_),
    .Y(_05178_),
    .A1(net3309),
    .A2(_05172_));
 sg13g2_o21ai_1 _11422_ (.B1(_05160_),
    .Y(_01353_),
    .A1(net3874),
    .A2(_05178_));
 sg13g2_nand2_1 _11423_ (.Y(_05179_),
    .A(\cpu.PCreg1[10] ),
    .B(net3873));
 sg13g2_and2_1 _11424_ (.A(_05151_),
    .B(_05164_),
    .X(_05180_));
 sg13g2_and2_1 _11425_ (.A(_05147_),
    .B(_05180_),
    .X(_05181_));
 sg13g2_o21ai_1 _11426_ (.B1(_05165_),
    .Y(_05182_),
    .A1(\cpu.PCci[9] ),
    .A2(_05162_));
 sg13g2_nand2_1 _11427_ (.Y(_05183_),
    .A(_05163_),
    .B(_05182_));
 sg13g2_a221oi_1 _11428_ (.B2(_05110_),
    .C1(_05183_),
    .B1(_05181_),
    .A1(_05146_),
    .Y(_05184_),
    .A2(_05180_));
 sg13g2_nand2_1 _11429_ (.Y(_05185_),
    .A(\cpu.Bimm[10] ),
    .B(net3415));
 sg13g2_o21ai_1 _11430_ (.B1(_05185_),
    .Y(_05186_),
    .A1(_00562_),
    .A2(net3114));
 sg13g2_xor2_1 _11431_ (.B(_05186_),
    .A(\cpu.PCci[10] ),
    .X(_05187_));
 sg13g2_nor2b_1 _11432_ (.A(_05184_),
    .B_N(_05187_),
    .Y(_05188_));
 sg13g2_nor2b_1 _11433_ (.A(_05187_),
    .B_N(_05184_),
    .Y(_05189_));
 sg13g2_or3_1 _11434_ (.A(net3112),
    .B(_05188_),
    .C(_05189_),
    .X(_05190_));
 sg13g2_xor2_1 _11435_ (.B(_05169_),
    .A(\cpu.PC[10] ),
    .X(_05191_));
 sg13g2_a21oi_1 _11436_ (.A1(net3112),
    .A2(_05191_),
    .Y(_05192_),
    .B1(net3424));
 sg13g2_a22oi_1 _11437_ (.Y(_05193_),
    .B1(_05190_),
    .B2(_05192_),
    .A2(_04035_),
    .A1(net3424));
 sg13g2_inv_1 _11438_ (.Y(_05194_),
    .A(_05193_));
 sg13g2_nand2b_1 _11439_ (.Y(_05195_),
    .B(net3248),
    .A_N(\irqvect[3][8] ));
 sg13g2_o21ai_1 _11440_ (.B1(_05195_),
    .Y(_05196_),
    .A1(\irqvect[2][8] ),
    .A2(net3251));
 sg13g2_mux2_1 _11441_ (.A0(\irqvect[0][8] ),
    .A1(\irqvect[1][8] ),
    .S(net3250),
    .X(_05197_));
 sg13g2_a21oi_1 _11442_ (.A1(net3320),
    .A2(_05197_),
    .Y(_05198_),
    .B1(net3258));
 sg13g2_o21ai_1 _11443_ (.B1(_05198_),
    .Y(_05199_),
    .A1(net3320),
    .A2(_05196_));
 sg13g2_o21ai_1 _11444_ (.B1(_05199_),
    .Y(_05200_),
    .A1(net3309),
    .A2(_05193_));
 sg13g2_o21ai_1 _11445_ (.B1(_05179_),
    .Y(_01354_),
    .A1(net3873),
    .A2(_05200_));
 sg13g2_nand2_1 _11446_ (.Y(_05201_),
    .A(net3645),
    .B(net3414));
 sg13g2_o21ai_1 _11447_ (.B1(_05201_),
    .Y(_05202_),
    .A1(_01690_),
    .A2(net3116));
 sg13g2_nor2_1 _11448_ (.A(\cpu.PCci[11] ),
    .B(_05202_),
    .Y(_05203_));
 sg13g2_xor2_1 _11449_ (.B(_05202_),
    .A(\cpu.PCci[11] ),
    .X(_05204_));
 sg13g2_a21o_1 _11450_ (.A2(_05186_),
    .A1(_01727_),
    .B1(_05188_),
    .X(_05205_));
 sg13g2_a21oi_1 _11451_ (.A1(\cpu.PC[10] ),
    .A2(_05169_),
    .Y(_05206_),
    .B1(\cpu.PC[11] ));
 sg13g2_and3_1 _11452_ (.X(_05207_),
    .A(\cpu.PC[11] ),
    .B(\cpu.PC[10] ),
    .C(_05169_));
 sg13g2_nor3_1 _11453_ (.A(net3107),
    .B(_05206_),
    .C(_05207_),
    .Y(_05208_));
 sg13g2_o21ai_1 _11454_ (.B1(net3107),
    .Y(_05209_),
    .A1(_05204_),
    .A2(_05205_));
 sg13g2_a21oi_1 _11455_ (.A1(_05204_),
    .A2(_05205_),
    .Y(_05210_),
    .B1(_05209_));
 sg13g2_o21ai_1 _11456_ (.B1(net3388),
    .Y(_05211_),
    .A1(_05208_),
    .A2(_05210_));
 sg13g2_nand2_1 _11457_ (.Y(_05212_),
    .A(net3422),
    .B(_04001_));
 sg13g2_and2_1 _11458_ (.A(_05211_),
    .B(_05212_),
    .X(_05213_));
 sg13g2_mux4_1 _11459_ (.S0(net3325),
    .A0(\irqvect[0][9] ),
    .A1(\irqvect[2][9] ),
    .A2(\irqvect[1][9] ),
    .A3(\irqvect[3][9] ),
    .S1(net3245),
    .X(_05214_));
 sg13g2_o21ai_1 _11460_ (.B1(net3707),
    .Y(_05215_),
    .A1(net3256),
    .A2(_05214_));
 sg13g2_a21oi_1 _11461_ (.A1(net3257),
    .A2(_05213_),
    .Y(_05216_),
    .B1(_05215_));
 sg13g2_a21o_1 _11462_ (.A2(net3873),
    .A1(\cpu.PCreg1[11] ),
    .B1(_05216_),
    .X(_01355_));
 sg13g2_a22oi_1 _11463_ (.Y(_05217_),
    .B1(_05202_),
    .B2(\cpu.PCci[11] ),
    .A2(_05186_),
    .A1(_01727_));
 sg13g2_nor2_1 _11464_ (.A(_05203_),
    .B(_05217_),
    .Y(_05218_));
 sg13g2_nand2_1 _11465_ (.Y(_05219_),
    .A(_05187_),
    .B(_05204_));
 sg13g2_nor2_1 _11466_ (.A(_05184_),
    .B(_05219_),
    .Y(_05220_));
 sg13g2_nor2_2 _11467_ (.A(net3640),
    .B(net3114),
    .Y(_05221_));
 sg13g2_nand2b_1 _11468_ (.Y(_05222_),
    .B(net3628),
    .A_N(net3114));
 sg13g2_nand2_1 _11469_ (.Y(_05223_),
    .A(net3699),
    .B(net3415));
 sg13g2_and2_1 _11470_ (.A(_05222_),
    .B(_05223_),
    .X(_05224_));
 sg13g2_o21ai_1 _11471_ (.B1(_05223_),
    .Y(_05225_),
    .A1(net3640),
    .A2(net3116));
 sg13g2_xor2_1 _11472_ (.B(_05225_),
    .A(\cpu.PCci[12] ),
    .X(_05226_));
 sg13g2_xnor2_1 _11473_ (.Y(_05227_),
    .A(\cpu.PCci[12] ),
    .B(_05225_));
 sg13g2_o21ai_1 _11474_ (.B1(_05226_),
    .Y(_05228_),
    .A1(_05218_),
    .A2(_05220_));
 sg13g2_or3_1 _11475_ (.A(_05218_),
    .B(_05220_),
    .C(_05226_),
    .X(_05229_));
 sg13g2_nand3_1 _11476_ (.B(_05228_),
    .C(_05229_),
    .A(net3106),
    .Y(_05230_));
 sg13g2_and2_1 _11477_ (.A(\cpu.PC[12] ),
    .B(_05207_),
    .X(_05231_));
 sg13g2_xor2_1 _11478_ (.B(_05207_),
    .A(\cpu.PC[12] ),
    .X(_05232_));
 sg13g2_a21oi_1 _11479_ (.A1(net3111),
    .A2(_05232_),
    .Y(_05233_),
    .B1(net3422));
 sg13g2_nand2_1 _11480_ (.Y(_05234_),
    .A(_05230_),
    .B(_05233_));
 sg13g2_o21ai_1 _11481_ (.B1(_05234_),
    .Y(_05235_),
    .A1(net3388),
    .A2(_04044_));
 sg13g2_mux2_1 _11482_ (.A0(\irqvect[0][10] ),
    .A1(\irqvect[1][10] ),
    .S(net3248),
    .X(_05236_));
 sg13g2_nand2_1 _11483_ (.Y(_05237_),
    .A(net3319),
    .B(_05236_));
 sg13g2_mux2_1 _11484_ (.A0(\irqvect[2][10] ),
    .A1(\irqvect[3][10] ),
    .S(net3248),
    .X(_05238_));
 sg13g2_a21oi_1 _11485_ (.A1(net3324),
    .A2(_05238_),
    .Y(_05239_),
    .B1(net3254));
 sg13g2_a221oi_1 _11486_ (.B2(_05239_),
    .C1(net3875),
    .B1(_05237_),
    .A1(net3254),
    .Y(_05240_),
    .A2(_05235_));
 sg13g2_a21o_1 _11487_ (.A2(net3875),
    .A1(\cpu.PCreg1[12] ),
    .B1(_05240_),
    .X(_01356_));
 sg13g2_and2_1 _11488_ (.A(_01728_),
    .B(_05225_),
    .X(_05241_));
 sg13g2_o21ai_1 _11489_ (.B1(_05228_),
    .Y(_05242_),
    .A1(_00569_),
    .A2(_05224_));
 sg13g2_nand2_1 _11490_ (.Y(_05243_),
    .A(net3697),
    .B(net3413));
 sg13g2_o21ai_1 _11491_ (.B1(_05243_),
    .Y(_05244_),
    .A1(net3640),
    .A2(net3116));
 sg13g2_and2_1 _11492_ (.A(\cpu.PCci[13] ),
    .B(_05244_),
    .X(_05245_));
 sg13g2_or2_1 _11493_ (.X(_05246_),
    .B(_05244_),
    .A(\cpu.PCci[13] ));
 sg13g2_xnor2_1 _11494_ (.Y(_05247_),
    .A(\cpu.PCci[13] ),
    .B(_05244_));
 sg13g2_inv_1 _11495_ (.Y(_05248_),
    .A(_05247_));
 sg13g2_o21ai_1 _11496_ (.B1(net3106),
    .Y(_05249_),
    .A1(_05242_),
    .A2(_05248_));
 sg13g2_a21oi_1 _11497_ (.A1(_05242_),
    .A2(_05248_),
    .Y(_05250_),
    .B1(_05249_));
 sg13g2_xnor2_1 _11498_ (.Y(_05251_),
    .A(\cpu.PC[13] ),
    .B(_05231_));
 sg13g2_o21ai_1 _11499_ (.B1(net3388),
    .Y(_05252_),
    .A1(net3106),
    .A2(_05251_));
 sg13g2_nand2_1 _11500_ (.Y(_05253_),
    .A(net3425),
    .B(_04051_));
 sg13g2_o21ai_1 _11501_ (.B1(_05253_),
    .Y(_05254_),
    .A1(_05250_),
    .A2(_05252_));
 sg13g2_mux4_1 _11502_ (.S0(net3322),
    .A0(\irqvect[0][11] ),
    .A1(\irqvect[2][11] ),
    .A2(\irqvect[1][11] ),
    .A3(\irqvect[3][11] ),
    .S1(net3247),
    .X(_05255_));
 sg13g2_o21ai_1 _11503_ (.B1(net3705),
    .Y(_05256_),
    .A1(net3253),
    .A2(_05255_));
 sg13g2_a21oi_1 _11504_ (.A1(net3256),
    .A2(_05254_),
    .Y(_05257_),
    .B1(_05256_));
 sg13g2_a21o_1 _11505_ (.A2(net3872),
    .A1(\cpu.PCreg1[13] ),
    .B1(_05257_),
    .X(_01357_));
 sg13g2_nand2_1 _11506_ (.Y(_05258_),
    .A(net3694),
    .B(net3413));
 sg13g2_o21ai_1 _11507_ (.B1(_05258_),
    .Y(_05259_),
    .A1(net3640),
    .A2(net3114));
 sg13g2_and2_1 _11508_ (.A(\cpu.PCci[14] ),
    .B(_05259_),
    .X(_05260_));
 sg13g2_xor2_1 _11509_ (.B(_05259_),
    .A(\cpu.PCci[14] ),
    .X(_05261_));
 sg13g2_or4_1 _11510_ (.A(_05203_),
    .B(_05217_),
    .C(_05227_),
    .D(_05247_),
    .X(_05262_));
 sg13g2_a21oi_1 _11511_ (.A1(_05241_),
    .A2(_05246_),
    .Y(_05263_),
    .B1(_05245_));
 sg13g2_and2_1 _11512_ (.A(_05262_),
    .B(_05263_),
    .X(_05264_));
 sg13g2_nand4_1 _11513_ (.B(_05204_),
    .C(_05226_),
    .A(_05187_),
    .Y(_05265_),
    .D(_05248_));
 sg13g2_o21ai_1 _11514_ (.B1(_05264_),
    .Y(_05266_),
    .A1(_05184_),
    .A2(_05265_));
 sg13g2_o21ai_1 _11515_ (.B1(net3106),
    .Y(_05267_),
    .A1(_05261_),
    .A2(_05266_));
 sg13g2_a21o_1 _11516_ (.A2(_05266_),
    .A1(_05261_),
    .B1(_05267_),
    .X(_05268_));
 sg13g2_nand3_1 _11517_ (.B(\cpu.PC[13] ),
    .C(_05231_),
    .A(\cpu.PC[14] ),
    .Y(_05269_));
 sg13g2_a21o_1 _11518_ (.A2(_05231_),
    .A1(\cpu.PC[13] ),
    .B1(\cpu.PC[14] ),
    .X(_05270_));
 sg13g2_nand3_1 _11519_ (.B(_05269_),
    .C(_05270_),
    .A(net3111),
    .Y(_05271_));
 sg13g2_nand3_1 _11520_ (.B(_05268_),
    .C(_05271_),
    .A(net3388),
    .Y(_05272_));
 sg13g2_o21ai_1 _11521_ (.B1(_05272_),
    .Y(_05273_),
    .A1(net3388),
    .A2(_03991_));
 sg13g2_mux4_1 _11522_ (.S0(net3322),
    .A0(\irqvect[0][12] ),
    .A1(\irqvect[2][12] ),
    .A2(\irqvect[1][12] ),
    .A3(\irqvect[3][12] ),
    .S1(net3246),
    .X(_05274_));
 sg13g2_o21ai_1 _11523_ (.B1(net3708),
    .Y(_05275_),
    .A1(net3253),
    .A2(_05274_));
 sg13g2_a21oi_1 _11524_ (.A1(net3257),
    .A2(_05273_),
    .Y(_05276_),
    .B1(_05275_));
 sg13g2_a21o_1 _11525_ (.A2(net3875),
    .A1(\cpu.PCreg1[14] ),
    .B1(_05276_),
    .X(_01358_));
 sg13g2_nand2_1 _11526_ (.Y(_05277_),
    .A(\cpu.PCreg1[15] ),
    .B(net3873));
 sg13g2_nand2_1 _11527_ (.Y(_05278_),
    .A(net3680),
    .B(net3413));
 sg13g2_o21ai_1 _11528_ (.B1(_05278_),
    .Y(_05279_),
    .A1(net3639),
    .A2(net3114));
 sg13g2_nor2_1 _11529_ (.A(\cpu.PCci[15] ),
    .B(_05279_),
    .Y(_05280_));
 sg13g2_xor2_1 _11530_ (.B(_05279_),
    .A(\cpu.PCci[15] ),
    .X(_05281_));
 sg13g2_a21o_1 _11531_ (.A2(_05266_),
    .A1(_05261_),
    .B1(_05260_),
    .X(_05282_));
 sg13g2_a21oi_1 _11532_ (.A1(_05281_),
    .A2(_05282_),
    .Y(_05283_),
    .B1(net3111));
 sg13g2_o21ai_1 _11533_ (.B1(_05283_),
    .Y(_05284_),
    .A1(_05281_),
    .A2(_05282_));
 sg13g2_nor2b_1 _11534_ (.A(_05269_),
    .B_N(\cpu.PC[15] ),
    .Y(_05285_));
 sg13g2_xnor2_1 _11535_ (.Y(_05286_),
    .A(\cpu.PC[15] ),
    .B(_05269_));
 sg13g2_a21oi_1 _11536_ (.A1(net3111),
    .A2(_05286_),
    .Y(_05287_),
    .B1(net3422));
 sg13g2_a22oi_1 _11537_ (.Y(_05288_),
    .B1(_05284_),
    .B2(_05287_),
    .A2(_03990_),
    .A1(net3422));
 sg13g2_nand2b_1 _11538_ (.Y(_05289_),
    .B(net3251),
    .A_N(\irqvect[3][13] ));
 sg13g2_o21ai_1 _11539_ (.B1(_05289_),
    .Y(_05290_),
    .A1(\irqvect[2][13] ),
    .A2(net3251));
 sg13g2_mux2_1 _11540_ (.A0(\irqvect[0][13] ),
    .A1(\irqvect[1][13] ),
    .S(net3251),
    .X(_05291_));
 sg13g2_a21oi_1 _11541_ (.A1(net3319),
    .A2(_05291_),
    .Y(_05292_),
    .B1(net3257));
 sg13g2_o21ai_1 _11542_ (.B1(_05292_),
    .Y(_05293_),
    .A1(net3319),
    .A2(_05290_));
 sg13g2_o21ai_1 _11543_ (.B1(_05293_),
    .Y(_05294_),
    .A1(net3308),
    .A2(_05288_));
 sg13g2_o21ai_1 _11544_ (.B1(_05277_),
    .Y(_01359_),
    .A1(net3873),
    .A2(_05294_));
 sg13g2_nand2_1 _11545_ (.Y(_05295_),
    .A(\cpu.PCreg1[16] ),
    .B(net3873));
 sg13g2_nand2_1 _11546_ (.Y(_05296_),
    .A(net3662),
    .B(net3413));
 sg13g2_o21ai_1 _11547_ (.B1(_05296_),
    .Y(_05297_),
    .A1(net3639),
    .A2(net3114));
 sg13g2_nand2_1 _11548_ (.Y(_05298_),
    .A(\cpu.PCci[16] ),
    .B(_05297_));
 sg13g2_xor2_1 _11549_ (.B(_05297_),
    .A(\cpu.PCci[16] ),
    .X(_05299_));
 sg13g2_inv_1 _11550_ (.Y(_05300_),
    .A(_05299_));
 sg13g2_and3_1 _11551_ (.X(_05301_),
    .A(_05261_),
    .B(_05266_),
    .C(_05281_));
 sg13g2_a22oi_1 _11552_ (.Y(_05302_),
    .B1(_05279_),
    .B2(\cpu.PCci[15] ),
    .A2(_05259_),
    .A1(\cpu.PCci[14] ));
 sg13g2_or2_1 _11553_ (.X(_05303_),
    .B(_05302_),
    .A(_05280_));
 sg13g2_inv_1 _11554_ (.Y(_05304_),
    .A(_05303_));
 sg13g2_nor3_1 _11555_ (.A(_05299_),
    .B(_05301_),
    .C(_05304_),
    .Y(_05305_));
 sg13g2_nor2_1 _11556_ (.A(net3111),
    .B(_05305_),
    .Y(_05306_));
 sg13g2_o21ai_1 _11557_ (.B1(_05299_),
    .Y(_05307_),
    .A1(_05301_),
    .A2(_05304_));
 sg13g2_nand2_1 _11558_ (.Y(_05308_),
    .A(\cpu.PC[16] ),
    .B(_05285_));
 sg13g2_xnor2_1 _11559_ (.Y(_05309_),
    .A(\cpu.PC[16] ),
    .B(_05285_));
 sg13g2_o21ai_1 _11560_ (.B1(net3388),
    .Y(_05310_),
    .A1(net3106),
    .A2(_05309_));
 sg13g2_a21oi_1 _11561_ (.A1(_05306_),
    .A2(_05307_),
    .Y(_05311_),
    .B1(_05310_));
 sg13g2_a21oi_2 _11562_ (.B1(_05311_),
    .Y(_05312_),
    .A2(_04032_),
    .A1(net3422));
 sg13g2_inv_1 _11563_ (.Y(_05313_),
    .A(_05312_));
 sg13g2_nand2b_1 _11564_ (.Y(_05314_),
    .B(net3248),
    .A_N(\irqvect[1][14] ));
 sg13g2_o21ai_1 _11565_ (.B1(_05314_),
    .Y(_05315_),
    .A1(\irqvect[0][14] ),
    .A2(net3248));
 sg13g2_mux2_1 _11566_ (.A0(\irqvect[2][14] ),
    .A1(\irqvect[3][14] ),
    .S(net3248),
    .X(_05316_));
 sg13g2_a21oi_1 _11567_ (.A1(net3323),
    .A2(_05316_),
    .Y(_05317_),
    .B1(net3254));
 sg13g2_o21ai_1 _11568_ (.B1(_05317_),
    .Y(_05318_),
    .A1(net3323),
    .A2(_05315_));
 sg13g2_o21ai_1 _11569_ (.B1(_05318_),
    .Y(_05319_),
    .A1(net3308),
    .A2(_05312_));
 sg13g2_o21ai_1 _11570_ (.B1(_05295_),
    .Y(_01360_),
    .A1(net3873),
    .A2(_05319_));
 sg13g2_nand2_1 _11571_ (.Y(_05320_),
    .A(\cpu.PCreg1[17] ),
    .B(net3873));
 sg13g2_nand2_1 _11572_ (.Y(_05321_),
    .A(net3655),
    .B(net3413));
 sg13g2_and2_1 _11573_ (.A(_05222_),
    .B(_05321_),
    .X(_05322_));
 sg13g2_o21ai_1 _11574_ (.B1(_05321_),
    .Y(_05323_),
    .A1(net3639),
    .A2(net3114));
 sg13g2_nor2_1 _11575_ (.A(_01731_),
    .B(_05322_),
    .Y(_05324_));
 sg13g2_xnor2_1 _11576_ (.Y(_05325_),
    .A(_01731_),
    .B(_05323_));
 sg13g2_xnor2_1 _11577_ (.Y(_05326_),
    .A(\cpu.PCci[17] ),
    .B(_05323_));
 sg13g2_nand3_1 _11578_ (.B(_05307_),
    .C(_05326_),
    .A(_05298_),
    .Y(_05327_));
 sg13g2_a21o_1 _11579_ (.A2(_05307_),
    .A1(_05298_),
    .B1(_05326_),
    .X(_05328_));
 sg13g2_nand3_1 _11580_ (.B(_05327_),
    .C(_05328_),
    .A(net3106),
    .Y(_05329_));
 sg13g2_nand3_1 _11581_ (.B(\cpu.PC[16] ),
    .C(_05285_),
    .A(\cpu.PC[17] ),
    .Y(_05330_));
 sg13g2_xnor2_1 _11582_ (.Y(_05331_),
    .A(\cpu.PC[17] ),
    .B(_05308_));
 sg13g2_a21oi_1 _11583_ (.A1(net3111),
    .A2(_05331_),
    .Y(_05332_),
    .B1(net3422));
 sg13g2_a22oi_1 _11584_ (.Y(_05333_),
    .B1(_05329_),
    .B2(_05332_),
    .A2(_04041_),
    .A1(net3422));
 sg13g2_nor2_1 _11585_ (.A(net3308),
    .B(_05333_),
    .Y(_05334_));
 sg13g2_mux4_1 _11586_ (.S0(net3322),
    .A0(\irqvect[0][15] ),
    .A1(\irqvect[2][15] ),
    .A2(\irqvect[1][15] ),
    .A3(\irqvect[3][15] ),
    .S1(net3247),
    .X(_05335_));
 sg13g2_o21ai_1 _11587_ (.B1(net3705),
    .Y(_05336_),
    .A1(net3254),
    .A2(_05335_));
 sg13g2_o21ai_1 _11588_ (.B1(_05320_),
    .Y(_01361_),
    .A1(_05334_),
    .A2(_05336_));
 sg13g2_nand2_1 _11589_ (.Y(_05337_),
    .A(\cpu.PCreg1[18] ),
    .B(net3872));
 sg13g2_and2_1 _11590_ (.A(\cpu.IR[18] ),
    .B(net3413),
    .X(_05338_));
 sg13g2_nor2_1 _11591_ (.A(_05221_),
    .B(_05338_),
    .Y(_05339_));
 sg13g2_o21ai_1 _11592_ (.B1(\cpu.PCci[18] ),
    .Y(_05340_),
    .A1(_05221_),
    .A2(_05338_));
 sg13g2_xnor2_1 _11593_ (.Y(_05341_),
    .A(\cpu.PCci[18] ),
    .B(_05339_));
 sg13g2_nand4_1 _11594_ (.B(_05281_),
    .C(_05299_),
    .A(_05261_),
    .Y(_05342_),
    .D(_05325_));
 sg13g2_or2_1 _11595_ (.X(_05343_),
    .B(_05342_),
    .A(_05265_));
 sg13g2_a21oi_1 _11596_ (.A1(_05262_),
    .A2(_05263_),
    .Y(_05344_),
    .B1(_05342_));
 sg13g2_a21oi_1 _11597_ (.A1(_01731_),
    .A2(_05322_),
    .Y(_05345_),
    .B1(_05298_));
 sg13g2_nor3_1 _11598_ (.A(_05300_),
    .B(_05303_),
    .C(_05326_),
    .Y(_05346_));
 sg13g2_nor4_1 _11599_ (.A(_05324_),
    .B(_05344_),
    .C(_05345_),
    .D(_05346_),
    .Y(_05347_));
 sg13g2_o21ai_1 _11600_ (.B1(_05347_),
    .Y(_05348_),
    .A1(_05184_),
    .A2(_05343_));
 sg13g2_xor2_1 _11601_ (.B(_05348_),
    .A(_05341_),
    .X(_05349_));
 sg13g2_nand2_1 _11602_ (.Y(_05350_),
    .A(net3105),
    .B(_05349_));
 sg13g2_nand2b_1 _11603_ (.Y(_05351_),
    .B(\cpu.PC[18] ),
    .A_N(_05330_));
 sg13g2_xnor2_1 _11604_ (.Y(_05352_),
    .A(\cpu.PC[18] ),
    .B(_05330_));
 sg13g2_a21oi_1 _11605_ (.A1(net3111),
    .A2(_05352_),
    .Y(_05353_),
    .B1(net3420));
 sg13g2_a22oi_1 _11606_ (.Y(_05354_),
    .B1(_05350_),
    .B2(_05353_),
    .A2(_03999_),
    .A1(net3420));
 sg13g2_inv_1 _11607_ (.Y(_05355_),
    .A(_05354_));
 sg13g2_nor2_1 _11608_ (.A(net3309),
    .B(_05354_),
    .Y(_05356_));
 sg13g2_mux4_1 _11609_ (.S0(net3322),
    .A0(\irqvect[0][16] ),
    .A1(\irqvect[2][16] ),
    .A2(\irqvect[1][16] ),
    .A3(\irqvect[3][16] ),
    .S1(net3247),
    .X(_05357_));
 sg13g2_o21ai_1 _11610_ (.B1(net3705),
    .Y(_05358_),
    .A1(net3254),
    .A2(_05357_));
 sg13g2_o21ai_1 _11611_ (.B1(_05337_),
    .Y(_01362_),
    .A1(_05356_),
    .A2(_05358_));
 sg13g2_nand2_1 _11612_ (.Y(_05359_),
    .A(net3420),
    .B(_04008_));
 sg13g2_nand2_1 _11613_ (.Y(_05360_),
    .A(\cpu.IR[19] ),
    .B(net3413));
 sg13g2_o21ai_1 _11614_ (.B1(_05360_),
    .Y(_05361_),
    .A1(net3639),
    .A2(net3114));
 sg13g2_xor2_1 _11615_ (.B(_05361_),
    .A(_00570_),
    .X(_05362_));
 sg13g2_nand2_1 _11616_ (.Y(_05363_),
    .A(_05340_),
    .B(_05362_));
 sg13g2_a21oi_1 _11617_ (.A1(_05341_),
    .A2(_05348_),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_nor2_1 _11618_ (.A(_05340_),
    .B(_05362_),
    .Y(_05365_));
 sg13g2_nor2b_1 _11619_ (.A(_05362_),
    .B_N(_05341_),
    .Y(_05366_));
 sg13g2_and2_1 _11620_ (.A(_05348_),
    .B(_05366_),
    .X(_05367_));
 sg13g2_nor4_1 _11621_ (.A(net3110),
    .B(_05364_),
    .C(_05365_),
    .D(_05367_),
    .Y(_05368_));
 sg13g2_nand2b_1 _11622_ (.Y(_05369_),
    .B(\cpu.PC[19] ),
    .A_N(_05351_));
 sg13g2_xor2_1 _11623_ (.B(_05351_),
    .A(\cpu.PC[19] ),
    .X(_05370_));
 sg13g2_o21ai_1 _11624_ (.B1(net3387),
    .Y(_05371_),
    .A1(net3105),
    .A2(_05370_));
 sg13g2_o21ai_1 _11625_ (.B1(_05359_),
    .Y(_05372_),
    .A1(_05368_),
    .A2(_05371_));
 sg13g2_mux4_1 _11626_ (.S0(net3321),
    .A0(\irqvect[0][17] ),
    .A1(\irqvect[2][17] ),
    .A2(\irqvect[1][17] ),
    .A3(\irqvect[3][17] ),
    .S1(net3245),
    .X(_05373_));
 sg13g2_o21ai_1 _11627_ (.B1(net3707),
    .Y(_05374_),
    .A1(net3255),
    .A2(_05373_));
 sg13g2_a21oi_1 _11628_ (.A1(net3255),
    .A2(_05372_),
    .Y(_05375_),
    .B1(_05374_));
 sg13g2_a21o_1 _11629_ (.A2(net3871),
    .A1(\cpu.PCreg1[19] ),
    .B1(_05375_),
    .X(_01363_));
 sg13g2_nand2_1 _11630_ (.Y(_05376_),
    .A(\cpu.PCreg1[20] ),
    .B(net3871));
 sg13g2_a21o_1 _11631_ (.A2(net3413),
    .A1(net3644),
    .B1(_05221_),
    .X(_05377_));
 sg13g2_nand2_1 _11632_ (.Y(_05378_),
    .A(\cpu.PCci[20] ),
    .B(net3102));
 sg13g2_inv_1 _11633_ (.Y(_05379_),
    .A(_05378_));
 sg13g2_xnor2_1 _11634_ (.Y(_05380_),
    .A(\cpu.PCci[20] ),
    .B(net3102));
 sg13g2_a21o_1 _11635_ (.A2(_05361_),
    .A1(\cpu.PCci[19] ),
    .B1(_05365_),
    .X(_05381_));
 sg13g2_a21oi_1 _11636_ (.A1(_05348_),
    .A2(_05366_),
    .Y(_05382_),
    .B1(_05381_));
 sg13g2_xor2_1 _11637_ (.B(_05382_),
    .A(_05380_),
    .X(_05383_));
 sg13g2_nand2_1 _11638_ (.Y(_05384_),
    .A(net3104),
    .B(_05383_));
 sg13g2_nand2b_1 _11639_ (.Y(_05385_),
    .B(\cpu.PC[20] ),
    .A_N(_05369_));
 sg13g2_xnor2_1 _11640_ (.Y(_05386_),
    .A(\cpu.PC[20] ),
    .B(_05369_));
 sg13g2_a21oi_1 _11641_ (.A1(net3109),
    .A2(_05386_),
    .Y(_05387_),
    .B1(net3418));
 sg13g2_a22oi_1 _11642_ (.Y(_05388_),
    .B1(_05384_),
    .B2(_05387_),
    .A2(_04004_),
    .A1(net3418));
 sg13g2_inv_1 _11643_ (.Y(_05389_),
    .A(_05388_));
 sg13g2_nor2_1 _11644_ (.A(net3308),
    .B(_05388_),
    .Y(_05390_));
 sg13g2_mux4_1 _11645_ (.S0(net3321),
    .A0(\irqvect[0][18] ),
    .A1(\irqvect[2][18] ),
    .A2(\irqvect[1][18] ),
    .A3(\irqvect[3][18] ),
    .S1(net3245),
    .X(_05391_));
 sg13g2_o21ai_1 _11646_ (.B1(net3705),
    .Y(_05392_),
    .A1(net3253),
    .A2(_05391_));
 sg13g2_o21ai_1 _11647_ (.B1(_05376_),
    .Y(_01364_),
    .A1(_05390_),
    .A2(_05392_));
 sg13g2_nand2_1 _11648_ (.Y(_05393_),
    .A(\cpu.PCreg1[21] ),
    .B(net3872));
 sg13g2_xnor2_1 _11649_ (.Y(_05394_),
    .A(\cpu.PCci[21] ),
    .B(net3103));
 sg13g2_o21ai_1 _11650_ (.B1(_05378_),
    .Y(_05395_),
    .A1(_05380_),
    .A2(_05382_));
 sg13g2_xnor2_1 _11651_ (.Y(_05396_),
    .A(_05394_),
    .B(_05395_));
 sg13g2_nand2_1 _11652_ (.Y(_05397_),
    .A(net3104),
    .B(_05396_));
 sg13g2_nor2b_1 _11653_ (.A(_05385_),
    .B_N(\cpu.PC[21] ),
    .Y(_05398_));
 sg13g2_xnor2_1 _11654_ (.Y(_05399_),
    .A(\cpu.PC[21] ),
    .B(_05385_));
 sg13g2_a21oi_1 _11655_ (.A1(net3109),
    .A2(_05399_),
    .Y(_05400_),
    .B1(net3418));
 sg13g2_a22oi_1 _11656_ (.Y(_05401_),
    .B1(_05397_),
    .B2(_05400_),
    .A2(_04009_),
    .A1(net3418));
 sg13g2_nor2_1 _11657_ (.A(net3309),
    .B(_05401_),
    .Y(_05402_));
 sg13g2_mux4_1 _11658_ (.S0(net3322),
    .A0(\irqvect[0][19] ),
    .A1(\irqvect[2][19] ),
    .A2(\irqvect[1][19] ),
    .A3(\irqvect[3][19] ),
    .S1(net3247),
    .X(_05403_));
 sg13g2_o21ai_1 _11659_ (.B1(net3705),
    .Y(_05404_),
    .A1(net3253),
    .A2(_05403_));
 sg13g2_o21ai_1 _11660_ (.B1(_05393_),
    .Y(_01365_),
    .A1(_05402_),
    .A2(_05404_));
 sg13g2_nand2_1 _11661_ (.Y(_05405_),
    .A(\cpu.PCci[22] ),
    .B(net3102));
 sg13g2_xor2_1 _11662_ (.B(net3102),
    .A(\cpu.PCci[22] ),
    .X(_05406_));
 sg13g2_inv_1 _11663_ (.Y(_05407_),
    .A(_05406_));
 sg13g2_nor2_1 _11664_ (.A(_05380_),
    .B(_05394_),
    .Y(_05408_));
 sg13g2_a221oi_1 _11665_ (.B2(_05408_),
    .C1(_05379_),
    .B1(_05381_),
    .A1(\cpu.PCci[21] ),
    .Y(_05409_),
    .A2(net3103));
 sg13g2_and2_1 _11666_ (.A(_05366_),
    .B(_05408_),
    .X(_05410_));
 sg13g2_nand2_1 _11667_ (.Y(_05411_),
    .A(_05366_),
    .B(_05408_));
 sg13g2_a21oi_1 _11668_ (.A1(_05381_),
    .A2(_05408_),
    .Y(_05412_),
    .B1(_05379_));
 sg13g2_inv_1 _11669_ (.Y(_05413_),
    .A(_05412_));
 sg13g2_a221oi_1 _11670_ (.B2(_05348_),
    .C1(_05413_),
    .B1(_05410_),
    .A1(\cpu.PCci[21] ),
    .Y(_05414_),
    .A2(net3103));
 sg13g2_xnor2_1 _11671_ (.Y(_05415_),
    .A(_05407_),
    .B(_05414_));
 sg13g2_nand2_1 _11672_ (.Y(_05416_),
    .A(\cpu.PC[22] ),
    .B(_05398_));
 sg13g2_xor2_1 _11673_ (.B(_05398_),
    .A(\cpu.PC[22] ),
    .X(_05417_));
 sg13g2_a21oi_1 _11674_ (.A1(net3109),
    .A2(_05417_),
    .Y(_05418_),
    .B1(net3418));
 sg13g2_o21ai_1 _11675_ (.B1(_05418_),
    .Y(_05419_),
    .A1(net3109),
    .A2(_05415_));
 sg13g2_o21ai_1 _11676_ (.B1(_05419_),
    .Y(_05420_),
    .A1(net3387),
    .A2(_04012_));
 sg13g2_mux4_1 _11677_ (.S0(net3321),
    .A0(\irqvect[0][20] ),
    .A1(\irqvect[2][20] ),
    .A2(\irqvect[1][20] ),
    .A3(\irqvect[3][20] ),
    .S1(net3245),
    .X(_05421_));
 sg13g2_o21ai_1 _11678_ (.B1(net3705),
    .Y(_05422_),
    .A1(net3253),
    .A2(_05421_));
 sg13g2_a21oi_1 _11679_ (.A1(net3256),
    .A2(_05420_),
    .Y(_05423_),
    .B1(_05422_));
 sg13g2_a21o_1 _11680_ (.A2(net3871),
    .A1(\cpu.PCreg1[22] ),
    .B1(_05423_),
    .X(_01366_));
 sg13g2_and2_1 _11681_ (.A(_00571_),
    .B(net3102),
    .X(_05424_));
 sg13g2_xnor2_1 _11682_ (.Y(_05425_),
    .A(_00571_),
    .B(net3102));
 sg13g2_o21ai_1 _11683_ (.B1(_05405_),
    .Y(_05426_),
    .A1(_05407_),
    .A2(_05414_));
 sg13g2_o21ai_1 _11684_ (.B1(net3104),
    .Y(_05427_),
    .A1(_05425_),
    .A2(_05426_));
 sg13g2_a21oi_1 _11685_ (.A1(_05425_),
    .A2(_05426_),
    .Y(_05428_),
    .B1(_05427_));
 sg13g2_nor2b_1 _11686_ (.A(_05416_),
    .B_N(\cpu.PC[23] ),
    .Y(_05429_));
 sg13g2_xor2_1 _11687_ (.B(_05416_),
    .A(\cpu.PC[23] ),
    .X(_05430_));
 sg13g2_o21ai_1 _11688_ (.B1(net3387),
    .Y(_05431_),
    .A1(net3105),
    .A2(_05430_));
 sg13g2_nand2_1 _11689_ (.Y(_05432_),
    .A(net3419),
    .B(_03983_));
 sg13g2_o21ai_1 _11690_ (.B1(_05432_),
    .Y(_05433_),
    .A1(_05428_),
    .A2(_05431_));
 sg13g2_mux2_1 _11691_ (.A0(\irqvect[2][21] ),
    .A1(\irqvect[3][21] ),
    .S(net3246),
    .X(_05434_));
 sg13g2_mux2_1 _11692_ (.A0(\irqvect[0][21] ),
    .A1(\irqvect[1][21] ),
    .S(net3246),
    .X(_05435_));
 sg13g2_nand2_1 _11693_ (.Y(_05436_),
    .A(net3319),
    .B(_05435_));
 sg13g2_a21oi_1 _11694_ (.A1(net3321),
    .A2(_05434_),
    .Y(_05437_),
    .B1(net3255));
 sg13g2_a221oi_1 _11695_ (.B2(_05437_),
    .C1(net3871),
    .B1(_05436_),
    .A1(net3255),
    .Y(_05438_),
    .A2(_05433_));
 sg13g2_a21o_1 _11696_ (.A2(net3871),
    .A1(\cpu.PCreg1[23] ),
    .B1(_05438_),
    .X(_01367_));
 sg13g2_nand2_1 _11697_ (.Y(_05439_),
    .A(\cpu.PCreg1[24] ),
    .B(net3872));
 sg13g2_and2_1 _11698_ (.A(\cpu.PCci[24] ),
    .B(net3103),
    .X(_05440_));
 sg13g2_xor2_1 _11699_ (.B(net3103),
    .A(\cpu.PCci[24] ),
    .X(_05441_));
 sg13g2_a22oi_1 _11700_ (.Y(_05442_),
    .B1(_05424_),
    .B2(\cpu.PCci[22] ),
    .A2(net3102),
    .A1(\cpu.PCci[23] ));
 sg13g2_nand2_1 _11701_ (.Y(_05443_),
    .A(_05406_),
    .B(_05425_));
 sg13g2_o21ai_1 _11702_ (.B1(_05442_),
    .Y(_05444_),
    .A1(_05414_),
    .A2(_05443_));
 sg13g2_o21ai_1 _11703_ (.B1(net3104),
    .Y(_05445_),
    .A1(_05441_),
    .A2(_05444_));
 sg13g2_a21o_1 _11704_ (.A2(_05444_),
    .A1(_05441_),
    .B1(_05445_),
    .X(_05446_));
 sg13g2_and2_1 _11705_ (.A(\cpu.PC[24] ),
    .B(_05429_),
    .X(_05447_));
 sg13g2_xor2_1 _11706_ (.B(_05429_),
    .A(\cpu.PC[24] ),
    .X(_05448_));
 sg13g2_a21oi_1 _11707_ (.A1(net3109),
    .A2(_05448_),
    .Y(_05449_),
    .B1(net3418));
 sg13g2_a22oi_1 _11708_ (.Y(_05450_),
    .B1(_05446_),
    .B2(_05449_),
    .A2(_04039_),
    .A1(net3418));
 sg13g2_nor2_1 _11709_ (.A(net3309),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_mux4_1 _11710_ (.S0(net3321),
    .A0(\irqvect[0][22] ),
    .A1(\irqvect[2][22] ),
    .A2(\irqvect[1][22] ),
    .A3(\irqvect[3][22] ),
    .S1(net3245),
    .X(_05452_));
 sg13g2_o21ai_1 _11711_ (.B1(net3707),
    .Y(_05453_),
    .A1(net3255),
    .A2(_05452_));
 sg13g2_o21ai_1 _11712_ (.B1(_05439_),
    .Y(_01368_),
    .A1(_05451_),
    .A2(_05453_));
 sg13g2_xor2_1 _11713_ (.B(_05447_),
    .A(\cpu.PC[25] ),
    .X(_05454_));
 sg13g2_a21oi_1 _11714_ (.A1(net3109),
    .A2(_05454_),
    .Y(_05455_),
    .B1(net3419));
 sg13g2_a21oi_1 _11715_ (.A1(_05441_),
    .A2(_05444_),
    .Y(_05456_),
    .B1(_05440_));
 sg13g2_xor2_1 _11716_ (.B(net3103),
    .A(\cpu.PCci[25] ),
    .X(_05457_));
 sg13g2_xor2_1 _11717_ (.B(_05457_),
    .A(_05456_),
    .X(_05458_));
 sg13g2_o21ai_1 _11718_ (.B1(_05455_),
    .Y(_05459_),
    .A1(net3109),
    .A2(_05458_));
 sg13g2_nand2_1 _11719_ (.Y(_05460_),
    .A(net3418),
    .B(_04045_));
 sg13g2_a21oi_1 _11720_ (.A1(_05459_),
    .A2(_05460_),
    .Y(_05461_),
    .B1(net3308));
 sg13g2_mux4_1 _11721_ (.S0(net3321),
    .A0(\irqvect[0][23] ),
    .A1(\irqvect[2][23] ),
    .A2(\irqvect[1][23] ),
    .A3(\irqvect[3][23] ),
    .S1(net3245),
    .X(_05462_));
 sg13g2_o21ai_1 _11722_ (.B1(net3707),
    .Y(_05463_),
    .A1(net3255),
    .A2(_05462_));
 sg13g2_nand2_1 _11723_ (.Y(_05464_),
    .A(\cpu.PCreg1[25] ),
    .B(net3872));
 sg13g2_o21ai_1 _11724_ (.B1(_05464_),
    .Y(_01369_),
    .A1(_05461_),
    .A2(_05463_));
 sg13g2_nand4_1 _11725_ (.B(_05425_),
    .C(_05441_),
    .A(_05406_),
    .Y(_05465_),
    .D(_05457_));
 sg13g2_o21ai_1 _11726_ (.B1(net3102),
    .Y(_05466_),
    .A1(\cpu.PCci[24] ),
    .A2(\cpu.PCci[25] ));
 sg13g2_and2_1 _11727_ (.A(_05442_),
    .B(_05466_),
    .X(_05467_));
 sg13g2_o21ai_1 _11728_ (.B1(_05467_),
    .Y(_05468_),
    .A1(_05409_),
    .A2(_05465_));
 sg13g2_nor2_1 _11729_ (.A(_05411_),
    .B(_05465_),
    .Y(_05469_));
 sg13g2_a21oi_1 _11730_ (.A1(_05348_),
    .A2(_05469_),
    .Y(_05470_),
    .B1(_05468_));
 sg13g2_a21o_1 _11731_ (.A2(_05469_),
    .A1(_05348_),
    .B1(_05468_),
    .X(_05471_));
 sg13g2_and2_1 _11732_ (.A(\cpu.PCci[26] ),
    .B(net3100),
    .X(_05472_));
 sg13g2_xor2_1 _11733_ (.B(net3100),
    .A(\cpu.PCci[26] ),
    .X(_05473_));
 sg13g2_a21oi_1 _11734_ (.A1(_05471_),
    .A2(_05473_),
    .Y(_05474_),
    .B1(net3109));
 sg13g2_o21ai_1 _11735_ (.B1(_05474_),
    .Y(_05475_),
    .A1(_05471_),
    .A2(_05473_));
 sg13g2_a21oi_1 _11736_ (.A1(\cpu.PC[25] ),
    .A2(_05447_),
    .Y(_05476_),
    .B1(\cpu.PC[26] ));
 sg13g2_and3_1 _11737_ (.X(_05477_),
    .A(\cpu.PC[25] ),
    .B(\cpu.PC[26] ),
    .C(_05447_));
 sg13g2_or3_1 _11738_ (.A(net3105),
    .B(_05476_),
    .C(_05477_),
    .X(_05478_));
 sg13g2_a21oi_1 _11739_ (.A1(_05475_),
    .A2(_05478_),
    .Y(_05479_),
    .B1(net3419));
 sg13g2_a21oi_2 _11740_ (.B1(_05479_),
    .Y(_05480_),
    .A2(_03995_),
    .A1(net3419));
 sg13g2_mux4_1 _11741_ (.S0(net3321),
    .A0(\irqvect[0][24] ),
    .A1(\irqvect[2][24] ),
    .A2(\irqvect[1][24] ),
    .A3(\irqvect[3][24] ),
    .S1(net3245),
    .X(_05481_));
 sg13g2_o21ai_1 _11742_ (.B1(net3707),
    .Y(_05482_),
    .A1(net3255),
    .A2(_05481_));
 sg13g2_a21oi_1 _11743_ (.A1(net3256),
    .A2(_05480_),
    .Y(_05483_),
    .B1(_05482_));
 sg13g2_a21o_1 _11744_ (.A2(net3872),
    .A1(\cpu.PCreg1[26] ),
    .B1(_05483_),
    .X(_01370_));
 sg13g2_xnor2_1 _11745_ (.Y(_05484_),
    .A(\cpu.PC[27] ),
    .B(_05477_));
 sg13g2_nand2_1 _11746_ (.Y(_05485_),
    .A(net3110),
    .B(_05484_));
 sg13g2_a21oi_1 _11747_ (.A1(_05471_),
    .A2(_05473_),
    .Y(_05486_),
    .B1(_05472_));
 sg13g2_xor2_1 _11748_ (.B(net3101),
    .A(\cpu.PCci[27] ),
    .X(_05487_));
 sg13g2_xnor2_1 _11749_ (.Y(_05488_),
    .A(_05486_),
    .B(_05487_));
 sg13g2_o21ai_1 _11750_ (.B1(_05485_),
    .Y(_05489_),
    .A1(net3110),
    .A2(_05488_));
 sg13g2_mux2_2 _11751_ (.A0(_04011_),
    .A1(_05489_),
    .S(net3387),
    .X(_05490_));
 sg13g2_mux2_1 _11752_ (.A0(\irqvect[0][25] ),
    .A1(\irqvect[1][25] ),
    .S(net3251),
    .X(_05491_));
 sg13g2_a21oi_1 _11753_ (.A1(_01733_),
    .A2(_04079_),
    .Y(_05492_),
    .B1(net3320));
 sg13g2_o21ai_1 _11754_ (.B1(_05492_),
    .Y(_05493_),
    .A1(\irqvect[2][25] ),
    .A2(net3248));
 sg13g2_a21oi_1 _11755_ (.A1(net3319),
    .A2(_05491_),
    .Y(_05494_),
    .B1(net3254));
 sg13g2_a221oi_1 _11756_ (.B2(_05494_),
    .C1(net3875),
    .B1(_05493_),
    .A1(net3254),
    .Y(_05495_),
    .A2(_05490_));
 sg13g2_a21o_1 _11757_ (.A2(net3875),
    .A1(\cpu.PCreg1[27] ),
    .B1(_05495_),
    .X(_01371_));
 sg13g2_nor2_1 _11758_ (.A(net3387),
    .B(_04015_),
    .Y(_05496_));
 sg13g2_o21ai_1 _11759_ (.B1(net3100),
    .Y(_05497_),
    .A1(\cpu.PCci[26] ),
    .A2(\cpu.PCci[27] ));
 sg13g2_nand2_1 _11760_ (.Y(_05498_),
    .A(_05473_),
    .B(_05487_));
 sg13g2_o21ai_1 _11761_ (.B1(_05497_),
    .Y(_05499_),
    .A1(_05470_),
    .A2(_05498_));
 sg13g2_and2_1 _11762_ (.A(\cpu.PCci[28] ),
    .B(net3101),
    .X(_05500_));
 sg13g2_xor2_1 _11763_ (.B(net3101),
    .A(\cpu.PCci[28] ),
    .X(_05501_));
 sg13g2_xnor2_1 _11764_ (.Y(_05502_),
    .A(_05499_),
    .B(_05501_));
 sg13g2_nand3_1 _11765_ (.B(\cpu.PC[28] ),
    .C(_05477_),
    .A(\cpu.PC[27] ),
    .Y(_05503_));
 sg13g2_a21o_1 _11766_ (.A2(_05477_),
    .A1(\cpu.PC[27] ),
    .B1(\cpu.PC[28] ),
    .X(_05504_));
 sg13g2_a21oi_1 _11767_ (.A1(_05503_),
    .A2(_05504_),
    .Y(_05505_),
    .B1(net3104));
 sg13g2_a21oi_1 _11768_ (.A1(net3104),
    .A2(_05502_),
    .Y(_05506_),
    .B1(_05505_));
 sg13g2_a21oi_2 _11769_ (.B1(_05496_),
    .Y(_05507_),
    .A2(_05506_),
    .A1(net3387));
 sg13g2_mux4_1 _11770_ (.S0(net3321),
    .A0(\irqvect[0][26] ),
    .A1(\irqvect[2][26] ),
    .A2(\irqvect[1][26] ),
    .A3(\irqvect[3][26] ),
    .S1(net3245),
    .X(_05508_));
 sg13g2_o21ai_1 _11771_ (.B1(net3707),
    .Y(_05509_),
    .A1(net3255),
    .A2(_05508_));
 sg13g2_a21oi_1 _11772_ (.A1(net3256),
    .A2(_05507_),
    .Y(_05510_),
    .B1(_05509_));
 sg13g2_a21o_1 _11773_ (.A2(net3874),
    .A1(\cpu.PCreg1[28] ),
    .B1(_05510_),
    .X(_01372_));
 sg13g2_nor2b_1 _11774_ (.A(_05503_),
    .B_N(\cpu.PC[29] ),
    .Y(_05511_));
 sg13g2_xnor2_1 _11775_ (.Y(_05512_),
    .A(\cpu.PC[29] ),
    .B(_05503_));
 sg13g2_a21oi_1 _11776_ (.A1(net3110),
    .A2(_05512_),
    .Y(_05513_),
    .B1(net3421));
 sg13g2_a21oi_1 _11777_ (.A1(_05499_),
    .A2(_05501_),
    .Y(_05514_),
    .B1(_05500_));
 sg13g2_xor2_1 _11778_ (.B(net3100),
    .A(\cpu.PCci[29] ),
    .X(_05515_));
 sg13g2_xor2_1 _11779_ (.B(_05515_),
    .A(_05514_),
    .X(_05516_));
 sg13g2_o21ai_1 _11780_ (.B1(_05513_),
    .Y(_05517_),
    .A1(net3110),
    .A2(_05516_));
 sg13g2_nand2_1 _11781_ (.Y(_05518_),
    .A(net3422),
    .B(_04048_));
 sg13g2_a21oi_1 _11782_ (.A1(_05517_),
    .A2(_05518_),
    .Y(_05519_),
    .B1(net3308));
 sg13g2_nand2b_1 _11783_ (.Y(_05520_),
    .B(net3246),
    .A_N(\irqvect[3][27] ));
 sg13g2_o21ai_1 _11784_ (.B1(_05520_),
    .Y(_05521_),
    .A1(\irqvect[2][27] ),
    .A2(net3246));
 sg13g2_mux2_1 _11785_ (.A0(\irqvect[0][27] ),
    .A1(\irqvect[1][27] ),
    .S(net3246),
    .X(_05522_));
 sg13g2_a21oi_1 _11786_ (.A1(net3319),
    .A2(_05522_),
    .Y(_05523_),
    .B1(net3253));
 sg13g2_o21ai_1 _11787_ (.B1(_05523_),
    .Y(_05524_),
    .A1(net3319),
    .A2(_05521_));
 sg13g2_nand2_1 _11788_ (.Y(_05525_),
    .A(net3708),
    .B(_05524_));
 sg13g2_nand2_1 _11789_ (.Y(_05526_),
    .A(\cpu.PCreg1[29] ),
    .B(net3871));
 sg13g2_o21ai_1 _11790_ (.B1(_05526_),
    .Y(_01373_),
    .A1(_05519_),
    .A2(_05525_));
 sg13g2_nand2_1 _11791_ (.Y(_05527_),
    .A(\cpu.PCreg1[30] ),
    .B(net3872));
 sg13g2_nand2_1 _11792_ (.Y(_05528_),
    .A(\cpu.PCci[30] ),
    .B(net3100));
 sg13g2_nor2_1 _11793_ (.A(\cpu.PCci[30] ),
    .B(net3100),
    .Y(_05529_));
 sg13g2_xor2_1 _11794_ (.B(net3100),
    .A(\cpu.PCci[30] ),
    .X(_05530_));
 sg13g2_nand2_1 _11795_ (.Y(_05531_),
    .A(_05501_),
    .B(_05515_));
 sg13g2_nor2_1 _11796_ (.A(_05498_),
    .B(_05531_),
    .Y(_05532_));
 sg13g2_o21ai_1 _11797_ (.B1(net3101),
    .Y(_05533_),
    .A1(\cpu.PCci[28] ),
    .A2(\cpu.PCci[29] ));
 sg13g2_o21ai_1 _11798_ (.B1(_05533_),
    .Y(_05534_),
    .A1(_05497_),
    .A2(_05531_));
 sg13g2_a21oi_1 _11799_ (.A1(_05471_),
    .A2(_05532_),
    .Y(_05535_),
    .B1(_05534_));
 sg13g2_xnor2_1 _11800_ (.Y(_05536_),
    .A(_05530_),
    .B(_05535_));
 sg13g2_nand2_1 _11801_ (.Y(_05537_),
    .A(\cpu.PC[30] ),
    .B(_05511_));
 sg13g2_xnor2_1 _11802_ (.Y(_05538_),
    .A(\cpu.PC[30] ),
    .B(_05511_));
 sg13g2_o21ai_1 _11803_ (.B1(net3387),
    .Y(_05539_),
    .A1(net3104),
    .A2(_05538_));
 sg13g2_a21oi_1 _11804_ (.A1(net3104),
    .A2(_05536_),
    .Y(_05540_),
    .B1(_05539_));
 sg13g2_nor2_1 _11805_ (.A(net3387),
    .B(_04014_),
    .Y(_05541_));
 sg13g2_nor2_1 _11806_ (.A(_05540_),
    .B(_05541_),
    .Y(_05542_));
 sg13g2_nand2b_1 _11807_ (.Y(_05543_),
    .B(net3247),
    .A_N(\irqvect[1][28] ));
 sg13g2_o21ai_1 _11808_ (.B1(_05543_),
    .Y(_05544_),
    .A1(\irqvect[0][28] ),
    .A2(net3247));
 sg13g2_mux2_1 _11809_ (.A0(\irqvect[2][28] ),
    .A1(\irqvect[3][28] ),
    .S(net3247),
    .X(_05545_));
 sg13g2_a21oi_1 _11810_ (.A1(net3322),
    .A2(_05545_),
    .Y(_05546_),
    .B1(net3253));
 sg13g2_o21ai_1 _11811_ (.B1(_05546_),
    .Y(_05547_),
    .A1(net3322),
    .A2(_05544_));
 sg13g2_o21ai_1 _11812_ (.B1(_05547_),
    .Y(_05548_),
    .A1(net3308),
    .A2(_05542_));
 sg13g2_o21ai_1 _11813_ (.B1(_05527_),
    .Y(_01374_),
    .A1(net3871),
    .A2(_05548_));
 sg13g2_nand2_2 _11814_ (.Y(_05549_),
    .A(net3421),
    .B(_04013_));
 sg13g2_o21ai_1 _11815_ (.B1(_05528_),
    .Y(_05550_),
    .A1(_05529_),
    .A2(_05535_));
 sg13g2_xor2_1 _11816_ (.B(net3100),
    .A(\cpu.PCci[31] ),
    .X(_05551_));
 sg13g2_xnor2_1 _11817_ (.Y(_05552_),
    .A(_05550_),
    .B(_05551_));
 sg13g2_xnor2_1 _11818_ (.Y(_05553_),
    .A(\cpu.PC[31] ),
    .B(_05537_));
 sg13g2_a21oi_1 _11819_ (.A1(net3110),
    .A2(_05553_),
    .Y(_05554_),
    .B1(net3421));
 sg13g2_o21ai_1 _11820_ (.B1(_05554_),
    .Y(_05555_),
    .A1(net3110),
    .A2(_05552_));
 sg13g2_a21oi_1 _11821_ (.A1(_05549_),
    .A2(_05555_),
    .Y(_05556_),
    .B1(net3308));
 sg13g2_mux4_1 _11822_ (.S0(net3322),
    .A0(\irqvect[0][29] ),
    .A1(\irqvect[2][29] ),
    .A2(\irqvect[1][29] ),
    .A3(\irqvect[3][29] ),
    .S1(net3247),
    .X(_05557_));
 sg13g2_o21ai_1 _11823_ (.B1(net3705),
    .Y(_05558_),
    .A1(net3253),
    .A2(_05557_));
 sg13g2_nand2_1 _11824_ (.Y(_05559_),
    .A(\cpu.PCreg1[31] ),
    .B(net3871));
 sg13g2_o21ai_1 _11825_ (.B1(_05559_),
    .Y(_01375_),
    .A1(_05556_),
    .A2(_05558_));
 sg13g2_nand2_1 _11826_ (.Y(_05560_),
    .A(_04910_),
    .B(_04917_));
 sg13g2_mux2_1 _11827_ (.A0(net3046),
    .A1(\cpu.regs[4][0] ),
    .S(net3144),
    .X(_01376_));
 sg13g2_mux2_1 _11828_ (.A0(net3041),
    .A1(\cpu.regs[4][1] ),
    .S(net3144),
    .X(_01377_));
 sg13g2_mux2_1 _11829_ (.A0(net3040),
    .A1(\cpu.regs[4][2] ),
    .S(net3143),
    .X(_01378_));
 sg13g2_mux2_1 _11830_ (.A0(net3005),
    .A1(\cpu.regs[4][3] ),
    .S(net3147),
    .X(_01379_));
 sg13g2_mux2_1 _11831_ (.A0(net3003),
    .A1(\cpu.regs[4][4] ),
    .S(net3144),
    .X(_01380_));
 sg13g2_mux2_1 _11832_ (.A0(net3029),
    .A1(\cpu.regs[4][5] ),
    .S(net3146),
    .X(_01381_));
 sg13g2_mux2_1 _11833_ (.A0(net3037),
    .A1(\cpu.regs[4][6] ),
    .S(net3144),
    .X(_01382_));
 sg13g2_mux2_1 _11834_ (.A0(net3044),
    .A1(\cpu.regs[4][7] ),
    .S(net3146),
    .X(_01383_));
 sg13g2_mux2_1 _11835_ (.A0(net3027),
    .A1(\cpu.regs[4][8] ),
    .S(net3146),
    .X(_01384_));
 sg13g2_mux2_1 _11836_ (.A0(net3026),
    .A1(\cpu.regs[4][9] ),
    .S(net3146),
    .X(_01385_));
 sg13g2_mux2_1 _11837_ (.A0(net3023),
    .A1(\cpu.regs[4][10] ),
    .S(net3147),
    .X(_01386_));
 sg13g2_mux2_1 _11838_ (.A0(net3021),
    .A1(\cpu.regs[4][11] ),
    .S(net3147),
    .X(_01387_));
 sg13g2_mux2_1 _11839_ (.A0(net3002),
    .A1(\cpu.regs[4][12] ),
    .S(net3143),
    .X(_01388_));
 sg13g2_mux2_1 _11840_ (.A0(net3019),
    .A1(\cpu.regs[4][13] ),
    .S(net3143),
    .X(_01389_));
 sg13g2_nand2_1 _11841_ (.Y(_05561_),
    .A(\cpu.regs[4][14] ),
    .B(net3146));
 sg13g2_o21ai_1 _11842_ (.B1(_05561_),
    .Y(_01390_),
    .A1(net3035),
    .A2(net3146));
 sg13g2_nand2_1 _11843_ (.Y(_05562_),
    .A(\cpu.regs[4][15] ),
    .B(net3146));
 sg13g2_o21ai_1 _11844_ (.B1(_05562_),
    .Y(_01391_),
    .A1(net3033),
    .A2(net3146));
 sg13g2_mux2_1 _11845_ (.A0(net2999),
    .A1(\cpu.regs[4][16] ),
    .S(net3143),
    .X(_01392_));
 sg13g2_nand2_1 _11846_ (.Y(_05563_),
    .A(\cpu.regs[4][17] ),
    .B(net3147));
 sg13g2_o21ai_1 _11847_ (.B1(_05563_),
    .Y(_01393_),
    .A1(net2997),
    .A2(net3147));
 sg13g2_mux2_1 _11848_ (.A0(net2995),
    .A1(\cpu.regs[4][18] ),
    .S(net3145),
    .X(_01394_));
 sg13g2_nand2_1 _11849_ (.Y(_05564_),
    .A(\cpu.regs[4][19] ),
    .B(net3147));
 sg13g2_o21ai_1 _11850_ (.B1(_05564_),
    .Y(_01395_),
    .A1(net2993),
    .A2(net3147));
 sg13g2_mux2_1 _11851_ (.A0(net2992),
    .A1(\cpu.regs[4][20] ),
    .S(net3143),
    .X(_01396_));
 sg13g2_mux2_1 _11852_ (.A0(net2989),
    .A1(\cpu.regs[4][21] ),
    .S(net3148),
    .X(_01397_));
 sg13g2_mux2_1 _11853_ (.A0(net3018),
    .A1(\cpu.regs[4][22] ),
    .S(net3145),
    .X(_01398_));
 sg13g2_mux2_1 _11854_ (.A0(net3015),
    .A1(\cpu.regs[4][23] ),
    .S(net3145),
    .X(_01399_));
 sg13g2_mux2_1 _11855_ (.A0(net2988),
    .A1(\cpu.regs[4][24] ),
    .S(net3145),
    .X(_01400_));
 sg13g2_mux2_1 _11856_ (.A0(net2985),
    .A1(\cpu.regs[4][25] ),
    .S(net3145),
    .X(_01401_));
 sg13g2_mux2_1 _11857_ (.A0(net3013),
    .A1(\cpu.regs[4][26] ),
    .S(net3143),
    .X(_01402_));
 sg13g2_mux2_1 _11858_ (.A0(net3011),
    .A1(\cpu.regs[4][27] ),
    .S(net3145),
    .X(_01403_));
 sg13g2_mux2_1 _11859_ (.A0(net2984),
    .A1(\cpu.regs[4][28] ),
    .S(net3145),
    .X(_01404_));
 sg13g2_mux2_1 _11860_ (.A0(net2981),
    .A1(\cpu.regs[4][29] ),
    .S(net3145),
    .X(_01405_));
 sg13g2_mux2_1 _11861_ (.A0(net3009),
    .A1(\cpu.regs[4][30] ),
    .S(net3143),
    .X(_01406_));
 sg13g2_mux2_1 _11862_ (.A0(net3007),
    .A1(\cpu.regs[4][31] ),
    .S(net3143),
    .X(_01407_));
 sg13g2_nor3_2 _11863_ (.A(_04122_),
    .B(_04896_),
    .C(_04903_),
    .Y(_05565_));
 sg13g2_mux2_1 _11864_ (.A0(\cpu.regs[3][0] ),
    .A1(net3046),
    .S(net3230),
    .X(_01408_));
 sg13g2_mux2_1 _11865_ (.A0(\cpu.regs[3][1] ),
    .A1(net3041),
    .S(net3230),
    .X(_01409_));
 sg13g2_mux2_1 _11866_ (.A0(\cpu.regs[3][2] ),
    .A1(net3040),
    .S(net3230),
    .X(_01410_));
 sg13g2_mux2_1 _11867_ (.A0(\cpu.regs[3][3] ),
    .A1(net3005),
    .S(net3229),
    .X(_01411_));
 sg13g2_mux2_1 _11868_ (.A0(\cpu.regs[3][4] ),
    .A1(net3003),
    .S(net3230),
    .X(_01412_));
 sg13g2_mux2_1 _11869_ (.A0(\cpu.regs[3][5] ),
    .A1(net3029),
    .S(net3229),
    .X(_01413_));
 sg13g2_mux2_1 _11870_ (.A0(\cpu.regs[3][6] ),
    .A1(net3037),
    .S(net3230),
    .X(_01414_));
 sg13g2_mux2_1 _11871_ (.A0(\cpu.regs[3][7] ),
    .A1(net3044),
    .S(net3229),
    .X(_01415_));
 sg13g2_mux2_1 _11872_ (.A0(\cpu.regs[3][8] ),
    .A1(net3027),
    .S(net3229),
    .X(_01416_));
 sg13g2_mux2_1 _11873_ (.A0(\cpu.regs[3][9] ),
    .A1(net3025),
    .S(net3228),
    .X(_01417_));
 sg13g2_mux2_1 _11874_ (.A0(\cpu.regs[3][10] ),
    .A1(net3023),
    .S(net3229),
    .X(_01418_));
 sg13g2_mux2_1 _11875_ (.A0(\cpu.regs[3][11] ),
    .A1(net3021),
    .S(net3229),
    .X(_01419_));
 sg13g2_mux2_1 _11876_ (.A0(\cpu.regs[3][12] ),
    .A1(net3001),
    .S(net3227),
    .X(_01420_));
 sg13g2_mux2_1 _11877_ (.A0(\cpu.regs[3][13] ),
    .A1(net3019),
    .S(net3227),
    .X(_01421_));
 sg13g2_nor2_1 _11878_ (.A(\cpu.regs[3][14] ),
    .B(net3228),
    .Y(_05566_));
 sg13g2_a21oi_1 _11879_ (.A1(net3035),
    .A2(net3228),
    .Y(_01422_),
    .B1(_05566_));
 sg13g2_nor2_1 _11880_ (.A(\cpu.regs[3][15] ),
    .B(net3228),
    .Y(_05567_));
 sg13g2_a21oi_1 _11881_ (.A1(net3033),
    .A2(net3228),
    .Y(_01423_),
    .B1(_05567_));
 sg13g2_mux2_1 _11882_ (.A0(\cpu.regs[3][16] ),
    .A1(net2999),
    .S(net3230),
    .X(_01424_));
 sg13g2_nor2_1 _11883_ (.A(\cpu.regs[3][17] ),
    .B(net3228),
    .Y(_05568_));
 sg13g2_a21oi_1 _11884_ (.A1(net2997),
    .A2(net3228),
    .Y(_01425_),
    .B1(_05568_));
 sg13g2_mux2_1 _11885_ (.A0(\cpu.regs[3][18] ),
    .A1(net2995),
    .S(net3226),
    .X(_01426_));
 sg13g2_nor2_1 _11886_ (.A(\cpu.regs[3][19] ),
    .B(net3229),
    .Y(_05569_));
 sg13g2_a21oi_1 _11887_ (.A1(net2993),
    .A2(net3228),
    .Y(_01427_),
    .B1(_05569_));
 sg13g2_mux2_1 _11888_ (.A0(\cpu.regs[3][20] ),
    .A1(net2991),
    .S(net3227),
    .X(_01428_));
 sg13g2_mux2_1 _11889_ (.A0(\cpu.regs[3][21] ),
    .A1(net2989),
    .S(net3226),
    .X(_01429_));
 sg13g2_mux2_1 _11890_ (.A0(\cpu.regs[3][22] ),
    .A1(net3018),
    .S(net3226),
    .X(_01430_));
 sg13g2_mux2_1 _11891_ (.A0(\cpu.regs[3][23] ),
    .A1(net3015),
    .S(net3226),
    .X(_01431_));
 sg13g2_mux2_1 _11892_ (.A0(\cpu.regs[3][24] ),
    .A1(net2987),
    .S(net3227),
    .X(_01432_));
 sg13g2_mux2_1 _11893_ (.A0(\cpu.regs[3][25] ),
    .A1(net2985),
    .S(net3226),
    .X(_01433_));
 sg13g2_mux2_1 _11894_ (.A0(\cpu.regs[3][26] ),
    .A1(net3013),
    .S(net3227),
    .X(_01434_));
 sg13g2_mux2_1 _11895_ (.A0(\cpu.regs[3][27] ),
    .A1(net3011),
    .S(net3226),
    .X(_01435_));
 sg13g2_mux2_1 _11896_ (.A0(\cpu.regs[3][28] ),
    .A1(net2984),
    .S(net3226),
    .X(_01436_));
 sg13g2_mux2_1 _11897_ (.A0(\cpu.regs[3][29] ),
    .A1(net2981),
    .S(net3226),
    .X(_01437_));
 sg13g2_mux2_1 _11898_ (.A0(\cpu.regs[3][30] ),
    .A1(net3009),
    .S(net3227),
    .X(_01438_));
 sg13g2_mux2_1 _11899_ (.A0(\cpu.regs[3][31] ),
    .A1(net3007),
    .S(net3227),
    .X(_01439_));
 sg13g2_mux2_1 _11900_ (.A0(_03329_),
    .A1(net921),
    .S(net3727),
    .X(_01440_));
 sg13g2_mux2_1 _11901_ (.A0(_03325_),
    .A1(net910),
    .S(net3727),
    .X(_01441_));
 sg13g2_mux2_1 _11902_ (.A0(_03321_),
    .A1(net923),
    .S(net3727),
    .X(_01442_));
 sg13g2_mux2_1 _11903_ (.A0(_03317_),
    .A1(net905),
    .S(net3727),
    .X(_01443_));
 sg13g2_mux2_1 _11904_ (.A0(_03314_),
    .A1(net918),
    .S(net3726),
    .X(_01444_));
 sg13g2_nand2_1 _11905_ (.Y(_05570_),
    .A(net893),
    .B(net3726));
 sg13g2_o21ai_1 _11906_ (.B1(_05570_),
    .Y(_01445_),
    .A1(net3725),
    .A2(_03309_));
 sg13g2_mux2_1 _11907_ (.A0(_03302_),
    .A1(net925),
    .S(net3727),
    .X(_01446_));
 sg13g2_mux2_1 _11908_ (.A0(_03299_),
    .A1(net912),
    .S(net3727),
    .X(_01447_));
 sg13g2_nor2_2 _11909_ (.A(net3626),
    .B(net3315),
    .Y(_05571_));
 sg13g2_and2_2 _11910_ (.A(net3631),
    .B(net3315),
    .X(_05572_));
 sg13g2_a22oi_1 _11911_ (.Y(_05573_),
    .B1(net3240),
    .B2(_01926_),
    .A2(net3244),
    .A1(\cpu.PCreg0[2] ));
 sg13g2_o21ai_1 _11912_ (.B1(_05573_),
    .Y(_01448_),
    .A1(net3636),
    .A2(_05056_));
 sg13g2_a22oi_1 _11913_ (.Y(_05574_),
    .B1(net3240),
    .B2(_01905_),
    .A2(net3244),
    .A1(\cpu.PCreg0[3] ));
 sg13g2_o21ai_1 _11914_ (.B1(_05574_),
    .Y(_01449_),
    .A1(net3637),
    .A2(_05070_));
 sg13g2_a22oi_1 _11915_ (.Y(_05575_),
    .B1(_05572_),
    .B2(_01887_),
    .A2(_05571_),
    .A1(\cpu.PCreg0[4] ));
 sg13g2_o21ai_1 _11916_ (.B1(_05575_),
    .Y(_01450_),
    .A1(net3635),
    .A2(_05087_));
 sg13g2_a22oi_1 _11917_ (.Y(_05576_),
    .B1(net3240),
    .B2(_01871_),
    .A2(net3244),
    .A1(\cpu.PCreg0[5] ));
 sg13g2_o21ai_1 _11918_ (.B1(_05576_),
    .Y(_01451_),
    .A1(net3636),
    .A2(_05104_));
 sg13g2_a22oi_1 _11919_ (.Y(_05577_),
    .B1(net3240),
    .B2(_01994_),
    .A2(net3244),
    .A1(\cpu.PCreg0[6] ));
 sg13g2_o21ai_1 _11920_ (.B1(_05577_),
    .Y(_01452_),
    .A1(net3636),
    .A2(_05120_));
 sg13g2_a22oi_1 _11921_ (.Y(_05578_),
    .B1(net3240),
    .B2(_01855_),
    .A2(net3244),
    .A1(\cpu.PCreg0[7] ));
 sg13g2_o21ai_1 _11922_ (.B1(_05578_),
    .Y(_01453_),
    .A1(net3636),
    .A2(_05137_));
 sg13g2_a22oi_1 _11923_ (.Y(_05579_),
    .B1(net3240),
    .B2(_02014_),
    .A2(net3244),
    .A1(\cpu.PCreg0[8] ));
 sg13g2_o21ai_1 _11924_ (.B1(_05579_),
    .Y(_01454_),
    .A1(net3635),
    .A2(_05156_));
 sg13g2_nand2_1 _11925_ (.Y(_05580_),
    .A(net3627),
    .B(_05172_));
 sg13g2_a22oi_1 _11926_ (.Y(_05581_),
    .B1(net3240),
    .B2(_02033_),
    .A2(net3244),
    .A1(\cpu.PCreg0[9] ));
 sg13g2_nand2_1 _11927_ (.Y(_01455_),
    .A(_05580_),
    .B(_05581_));
 sg13g2_a22oi_1 _11928_ (.Y(_05582_),
    .B1(net3240),
    .B2(_02053_),
    .A2(net3244),
    .A1(\cpu.PCreg0[10] ));
 sg13g2_o21ai_1 _11929_ (.B1(_05582_),
    .Y(_01456_),
    .A1(net3635),
    .A2(_05194_));
 sg13g2_a22oi_1 _11930_ (.Y(_05583_),
    .B1(net3239),
    .B2(_01839_),
    .A2(net3243),
    .A1(\cpu.PCreg0[11] ));
 sg13g2_o21ai_1 _11931_ (.B1(_05583_),
    .Y(_01457_),
    .A1(net3630),
    .A2(_05213_));
 sg13g2_a22oi_1 _11932_ (.Y(_05584_),
    .B1(net3239),
    .B2(_02078_),
    .A2(net3243),
    .A1(\cpu.PCreg0[12] ));
 sg13g2_o21ai_1 _11933_ (.B1(_05584_),
    .Y(_01458_),
    .A1(net3629),
    .A2(_05235_));
 sg13g2_a22oi_1 _11934_ (.Y(_05585_),
    .B1(net3238),
    .B2(_02097_),
    .A2(net3242),
    .A1(\cpu.PCreg0[13] ));
 sg13g2_o21ai_1 _11935_ (.B1(_05585_),
    .Y(_01459_),
    .A1(net3629),
    .A2(_05254_));
 sg13g2_a22oi_1 _11936_ (.Y(_05586_),
    .B1(net3239),
    .B2(_01824_),
    .A2(net3243),
    .A1(\cpu.PCreg0[14] ));
 sg13g2_o21ai_1 _11937_ (.B1(_05586_),
    .Y(_01460_),
    .A1(net3630),
    .A2(_05273_));
 sg13g2_nand2_1 _11938_ (.Y(_05587_),
    .A(net3627),
    .B(_05288_));
 sg13g2_a22oi_1 _11939_ (.Y(_05588_),
    .B1(net3239),
    .B2(_01807_),
    .A2(net3243),
    .A1(\cpu.PCreg0[15] ));
 sg13g2_nand2_1 _11940_ (.Y(_01461_),
    .A(_05587_),
    .B(_05588_));
 sg13g2_a22oi_1 _11941_ (.Y(_05589_),
    .B1(net3239),
    .B2(_02118_),
    .A2(net3243),
    .A1(\cpu.PCreg0[16] ));
 sg13g2_o21ai_1 _11942_ (.B1(_05589_),
    .Y(_01462_),
    .A1(net3630),
    .A2(_05313_));
 sg13g2_nand2_1 _11943_ (.Y(_05590_),
    .A(net3627),
    .B(_05333_));
 sg13g2_a22oi_1 _11944_ (.Y(_05591_),
    .B1(net3239),
    .B2(_02222_),
    .A2(net3243),
    .A1(\cpu.PCreg0[17] ));
 sg13g2_nand2_1 _11945_ (.Y(_01463_),
    .A(_05590_),
    .B(_05591_));
 sg13g2_a22oi_1 _11946_ (.Y(_05592_),
    .B1(net3237),
    .B2(_02205_),
    .A2(net3241),
    .A1(\cpu.PCreg0[18] ));
 sg13g2_o21ai_1 _11947_ (.B1(_05592_),
    .Y(_01464_),
    .A1(net3634),
    .A2(_05355_));
 sg13g2_a22oi_1 _11948_ (.Y(_05593_),
    .B1(net3237),
    .B2(_02242_),
    .A2(net3241),
    .A1(\cpu.PCreg0[19] ));
 sg13g2_o21ai_1 _11949_ (.B1(_05593_),
    .Y(_01465_),
    .A1(net3633),
    .A2(_05372_));
 sg13g2_a22oi_1 _11950_ (.Y(_05594_),
    .B1(net3238),
    .B2(_02185_),
    .A2(net3242),
    .A1(\cpu.PCreg0[20] ));
 sg13g2_o21ai_1 _11951_ (.B1(_05594_),
    .Y(_01466_),
    .A1(net3631),
    .A2(_05389_));
 sg13g2_nand2_1 _11952_ (.Y(_05595_),
    .A(net3626),
    .B(_05401_));
 sg13g2_a22oi_1 _11953_ (.Y(_05596_),
    .B1(net3237),
    .B2(_02171_),
    .A2(net3241),
    .A1(\cpu.PCreg0[21] ));
 sg13g2_nand2_1 _11954_ (.Y(_01467_),
    .A(_05595_),
    .B(_05596_));
 sg13g2_a22oi_1 _11955_ (.Y(_05597_),
    .B1(net3237),
    .B2(_02134_),
    .A2(net3241),
    .A1(\cpu.PCreg0[22] ));
 sg13g2_o21ai_1 _11956_ (.B1(_05597_),
    .Y(_01468_),
    .A1(net3632),
    .A2(_05420_));
 sg13g2_a22oi_1 _11957_ (.Y(_05598_),
    .B1(net3237),
    .B2(_02152_),
    .A2(net3241),
    .A1(\cpu.PCreg0[23] ));
 sg13g2_o21ai_1 _11958_ (.B1(_05598_),
    .Y(_01469_),
    .A1(net3632),
    .A2(_05433_));
 sg13g2_nand2_1 _11959_ (.Y(_05599_),
    .A(net3626),
    .B(_05450_));
 sg13g2_nand2_1 _11960_ (.Y(_05600_),
    .A(\cpu.PCreg0[24] ),
    .B(net3241));
 sg13g2_nand2_1 _11961_ (.Y(_05601_),
    .A(_02297_),
    .B(net3237));
 sg13g2_nand3_1 _11962_ (.B(_05600_),
    .C(_05601_),
    .A(_05599_),
    .Y(_01470_));
 sg13g2_nand3_1 _11963_ (.B(_05459_),
    .C(_05460_),
    .A(net3626),
    .Y(_05602_));
 sg13g2_a22oi_1 _11964_ (.Y(_05603_),
    .B1(net3237),
    .B2(_02314_),
    .A2(net3241),
    .A1(\cpu.PCreg0[25] ));
 sg13g2_nand2_1 _11965_ (.Y(_01471_),
    .A(_05602_),
    .B(_05603_));
 sg13g2_a22oi_1 _11966_ (.Y(_05604_),
    .B1(net3237),
    .B2(_02282_),
    .A2(net3241),
    .A1(\cpu.PCreg0[26] ));
 sg13g2_o21ai_1 _11967_ (.B1(_05604_),
    .Y(_01472_),
    .A1(net3633),
    .A2(_05480_));
 sg13g2_a22oi_1 _11968_ (.Y(_05605_),
    .B1(net3238),
    .B2(_02268_),
    .A2(net3242),
    .A1(\cpu.PCreg0[27] ));
 sg13g2_o21ai_1 _11969_ (.B1(_05605_),
    .Y(_01473_),
    .A1(net3633),
    .A2(_05490_));
 sg13g2_a22oi_1 _11970_ (.Y(_05606_),
    .B1(net3238),
    .B2(_02339_),
    .A2(net3242),
    .A1(\cpu.PCreg0[28] ));
 sg13g2_o21ai_1 _11971_ (.B1(_05606_),
    .Y(_01474_),
    .A1(net3633),
    .A2(_05507_));
 sg13g2_nand3_1 _11972_ (.B(_05517_),
    .C(_05518_),
    .A(net3626),
    .Y(_05607_));
 sg13g2_a22oi_1 _11973_ (.Y(_05608_),
    .B1(net3238),
    .B2(_02358_),
    .A2(net3242),
    .A1(\cpu.PCreg0[29] ));
 sg13g2_nand2_1 _11974_ (.Y(_01475_),
    .A(_05607_),
    .B(_05608_));
 sg13g2_nand2_1 _11975_ (.Y(_05609_),
    .A(net3626),
    .B(_05542_));
 sg13g2_a22oi_1 _11976_ (.Y(_05610_),
    .B1(net3238),
    .B2(_01791_),
    .A2(net3242),
    .A1(\cpu.PCreg0[30] ));
 sg13g2_nand2_1 _11977_ (.Y(_01476_),
    .A(_05609_),
    .B(_05610_));
 sg13g2_nand3_1 _11978_ (.B(_05549_),
    .C(_05555_),
    .A(net3626),
    .Y(_05611_));
 sg13g2_a22oi_1 _11979_ (.Y(_05612_),
    .B1(net3238),
    .B2(_02383_),
    .A2(net3242),
    .A1(\cpu.PCreg0[31] ));
 sg13g2_nand2_1 _11980_ (.Y(_01477_),
    .A(_05611_),
    .B(_05612_));
 sg13g2_nor3_2 _11981_ (.A(net3125),
    .B(_03445_),
    .C(_04868_),
    .Y(_05613_));
 sg13g2_mux2_1 _11982_ (.A0(\irqvect[3][0] ),
    .A1(net3326),
    .S(net3058),
    .X(_01478_));
 sg13g2_mux2_1 _11983_ (.A0(\irqvect[3][1] ),
    .A1(net3327),
    .S(net3060),
    .X(_01479_));
 sg13g2_nor2_1 _11984_ (.A(\irqvect[3][2] ),
    .B(net3059),
    .Y(_05614_));
 sg13g2_a21oi_1 _11985_ (.A1(_02928_),
    .A2(net3059),
    .Y(_01480_),
    .B1(_05614_));
 sg13g2_mux2_1 _11986_ (.A0(\irqvect[3][3] ),
    .A1(net3328),
    .S(net3060),
    .X(_01481_));
 sg13g2_mux2_1 _11987_ (.A0(\irqvect[3][4] ),
    .A1(net3329),
    .S(net3059),
    .X(_01482_));
 sg13g2_mux2_1 _11988_ (.A0(\irqvect[3][5] ),
    .A1(net3330),
    .S(net3060),
    .X(_01483_));
 sg13g2_nor2_1 _11989_ (.A(\irqvect[3][6] ),
    .B(net3059),
    .Y(_05615_));
 sg13g2_a21oi_1 _11990_ (.A1(_03267_),
    .A2(net3059),
    .Y(_01484_),
    .B1(_05615_));
 sg13g2_nor2_1 _11991_ (.A(\irqvect[3][7] ),
    .B(net3059),
    .Y(_05616_));
 sg13g2_a21oi_1 _11992_ (.A1(_03193_),
    .A2(net3059),
    .Y(_01485_),
    .B1(_05616_));
 sg13g2_nor2_1 _11993_ (.A(\irqvect[3][8] ),
    .B(net3060),
    .Y(_05617_));
 sg13g2_a21oi_1 _11994_ (.A1(_03120_),
    .A2(net3058),
    .Y(_01486_),
    .B1(_05617_));
 sg13g2_nor2_1 _11995_ (.A(\irqvect[3][9] ),
    .B(net3057),
    .Y(_05618_));
 sg13g2_a21oi_1 _11996_ (.A1(_03033_),
    .A2(net3057),
    .Y(_01487_),
    .B1(_05618_));
 sg13g2_nor2_1 _11997_ (.A(\irqvect[3][10] ),
    .B(net3058),
    .Y(_05619_));
 sg13g2_a21oi_1 _11998_ (.A1(_02947_),
    .A2(net3058),
    .Y(_01488_),
    .B1(_05619_));
 sg13g2_nor2_1 _11999_ (.A(\irqvect[3][11] ),
    .B(net3052),
    .Y(_05620_));
 sg13g2_a21oi_1 _12000_ (.A1(_02861_),
    .A2(net3052),
    .Y(_01489_),
    .B1(_05620_));
 sg13g2_nor2_1 _12001_ (.A(\irqvect[3][12] ),
    .B(net3056),
    .Y(_05621_));
 sg13g2_a21oi_1 _12002_ (.A1(_02778_),
    .A2(net3056),
    .Y(_01490_),
    .B1(_05621_));
 sg13g2_nor2_1 _12003_ (.A(\irqvect[3][13] ),
    .B(net3060),
    .Y(_05622_));
 sg13g2_a21oi_1 _12004_ (.A1(_02682_),
    .A2(net3060),
    .Y(_01491_),
    .B1(_05622_));
 sg13g2_nor2_1 _12005_ (.A(\irqvect[3][14] ),
    .B(net3058),
    .Y(_05623_));
 sg13g2_a21oi_1 _12006_ (.A1(_03288_),
    .A2(net3058),
    .Y(_01492_),
    .B1(_05623_));
 sg13g2_nor2_1 _12007_ (.A(\irqvect[3][15] ),
    .B(net3052),
    .Y(_05624_));
 sg13g2_a21oi_1 _12008_ (.A1(_03216_),
    .A2(net3052),
    .Y(_01493_),
    .B1(_05624_));
 sg13g2_nor2_1 _12009_ (.A(\irqvect[3][16] ),
    .B(net3052),
    .Y(_05625_));
 sg13g2_a21oi_1 _12010_ (.A1(_03142_),
    .A2(net3052),
    .Y(_01494_),
    .B1(_05625_));
 sg13g2_nor2_1 _12011_ (.A(\irqvect[3][17] ),
    .B(net3055),
    .Y(_05626_));
 sg13g2_a21oi_1 _12012_ (.A1(_03054_),
    .A2(net3054),
    .Y(_01495_),
    .B1(_05626_));
 sg13g2_nor2_1 _12013_ (.A(\irqvect[3][18] ),
    .B(net3054),
    .Y(_05627_));
 sg13g2_a21oi_1 _12014_ (.A1(_02967_),
    .A2(net3054),
    .Y(_01496_),
    .B1(_05627_));
 sg13g2_nor2_1 _12015_ (.A(\irqvect[3][19] ),
    .B(net3053),
    .Y(_05628_));
 sg13g2_a21oi_1 _12016_ (.A1(_02881_),
    .A2(net3053),
    .Y(_01497_),
    .B1(_05628_));
 sg13g2_nor2_1 _12017_ (.A(\irqvect[3][20] ),
    .B(net3054),
    .Y(_05629_));
 sg13g2_a21oi_1 _12018_ (.A1(_02798_),
    .A2(net3054),
    .Y(_01498_),
    .B1(_05629_));
 sg13g2_nor2_1 _12019_ (.A(\irqvect[3][21] ),
    .B(net3056),
    .Y(_05630_));
 sg13g2_a21oi_1 _12020_ (.A1(_02703_),
    .A2(net3056),
    .Y(_01499_),
    .B1(_05630_));
 sg13g2_nor2_1 _12021_ (.A(\irqvect[3][22] ),
    .B(net3055),
    .Y(_05631_));
 sg13g2_a21oi_1 _12022_ (.A1(_03269_),
    .A2(net3054),
    .Y(_01500_),
    .B1(_05631_));
 sg13g2_nor2_1 _12023_ (.A(\irqvect[3][23] ),
    .B(net3055),
    .Y(_05632_));
 sg13g2_a21oi_1 _12024_ (.A1(_03195_),
    .A2(net3055),
    .Y(_01501_),
    .B1(_05632_));
 sg13g2_nor2_1 _12025_ (.A(\irqvect[3][24] ),
    .B(net3055),
    .Y(_05633_));
 sg13g2_a21oi_1 _12026_ (.A1(_03122_),
    .A2(net3055),
    .Y(_01502_),
    .B1(_05633_));
 sg13g2_nor2_1 _12027_ (.A(\irqvect[3][25] ),
    .B(net3058),
    .Y(_05634_));
 sg13g2_a21oi_1 _12028_ (.A1(_03035_),
    .A2(net3058),
    .Y(_01503_),
    .B1(_05634_));
 sg13g2_nor2_1 _12029_ (.A(\irqvect[3][26] ),
    .B(net3054),
    .Y(_05635_));
 sg13g2_a21oi_1 _12030_ (.A1(_02949_),
    .A2(net3054),
    .Y(_01504_),
    .B1(_05635_));
 sg13g2_nor2_1 _12031_ (.A(\irqvect[3][27] ),
    .B(net3056),
    .Y(_05636_));
 sg13g2_a21oi_1 _12032_ (.A1(_02863_),
    .A2(net3056),
    .Y(_01505_),
    .B1(_05636_));
 sg13g2_nor2_1 _12033_ (.A(\irqvect[3][28] ),
    .B(net3052),
    .Y(_05637_));
 sg13g2_a21oi_1 _12034_ (.A1(_02780_),
    .A2(net3052),
    .Y(_01506_),
    .B1(_05637_));
 sg13g2_nor2_1 _12035_ (.A(\irqvect[3][29] ),
    .B(net3053),
    .Y(_05638_));
 sg13g2_a21oi_1 _12036_ (.A1(_02684_),
    .A2(net3053),
    .Y(_01507_),
    .B1(_05638_));
 sg13g2_inv_1 _12037_ (.Y(_00592_),
    .A(net3941));
 sg13g2_inv_1 _12038_ (.Y(_00593_),
    .A(net3941));
 sg13g2_inv_1 _12039_ (.Y(_00594_),
    .A(net3941));
 sg13g2_inv_1 _12040_ (.Y(_00595_),
    .A(net3942));
 sg13g2_inv_1 _12041_ (.Y(_00596_),
    .A(net3941));
 sg13g2_inv_1 _12042_ (.Y(_00597_),
    .A(net3940));
 sg13g2_inv_1 _12043_ (.Y(_00598_),
    .A(net3940));
 sg13g2_inv_1 _12044_ (.Y(_00599_),
    .A(net3938));
 sg13g2_inv_1 _12045_ (.Y(_00600_),
    .A(net3938));
 sg13g2_inv_1 _12046_ (.Y(_00601_),
    .A(net3938));
 sg13g2_inv_1 _12047_ (.Y(_00602_),
    .A(net3936));
 sg13g2_inv_1 _12048_ (.Y(_00603_),
    .A(net3936));
 sg13g2_inv_1 _12049_ (.Y(_00604_),
    .A(net3935));
 sg13g2_inv_1 _12050_ (.Y(_00605_),
    .A(net3935));
 sg13g2_inv_1 _12051_ (.Y(_00606_),
    .A(net3935));
 sg13g2_inv_1 _12052_ (.Y(_00607_),
    .A(net3937));
 sg13g2_inv_1 _12053_ (.Y(_00608_),
    .A(net3937));
 sg13g2_inv_1 _12054_ (.Y(_00609_),
    .A(net3939));
 sg13g2_inv_1 _12055_ (.Y(_00610_),
    .A(net3937));
 sg13g2_inv_1 _12056_ (.Y(_00611_),
    .A(net3937));
 sg13g2_inv_1 _12057_ (.Y(_00612_),
    .A(net3937));
 sg13g2_inv_1 _12058_ (.Y(_00613_),
    .A(net3937));
 sg13g2_inv_1 _12059_ (.Y(_00614_),
    .A(net3935));
 sg13g2_inv_1 _12060_ (.Y(_00615_),
    .A(net3935));
 sg13g2_inv_1 _12061_ (.Y(_00616_),
    .A(net3935));
 sg13g2_inv_1 _12062_ (.Y(_00617_),
    .A(net3935));
 sg13g2_inv_1 _12063_ (.Y(_00618_),
    .A(net3935));
 sg13g2_inv_1 _12064_ (.Y(_00619_),
    .A(net3936));
 sg13g2_inv_1 _12065_ (.Y(_00620_),
    .A(net3936));
 sg13g2_inv_1 _12066_ (.Y(_00621_),
    .A(net3936));
 sg13g2_inv_1 _12067_ (.Y(_00622_),
    .A(net3938));
 sg13g2_inv_1 _12068_ (.Y(_00623_),
    .A(net3938));
 sg13g2_inv_1 _12069_ (.Y(_00624_),
    .A(net3936));
 sg13g2_inv_1 _12070_ (.Y(_00625_),
    .A(net3936));
 sg13g2_inv_1 _12071_ (.Y(_00626_),
    .A(net3936));
 sg13g2_inv_1 _12072_ (.Y(_00627_),
    .A(net3938));
 sg13g2_inv_1 _12073_ (.Y(_00628_),
    .A(net3938));
 sg13g2_inv_1 _12074_ (.Y(_00629_),
    .A(net3938));
 sg13g2_inv_1 _12075_ (.Y(_00630_),
    .A(net3939));
 sg13g2_inv_1 _12076_ (.Y(_00631_),
    .A(net3940));
 sg13g2_inv_1 _12077_ (.Y(_00632_),
    .A(net3940));
 sg13g2_inv_1 _12078_ (.Y(_00633_),
    .A(net3944));
 sg13g2_inv_1 _12079_ (.Y(_00634_),
    .A(net3947));
 sg13g2_inv_1 _12080_ (.Y(_00635_),
    .A(net3946));
 sg13g2_inv_1 _12081_ (.Y(_00636_),
    .A(net3948));
 sg13g2_inv_1 _12082_ (.Y(_00637_),
    .A(net3949));
 sg13g2_inv_1 _12083_ (.Y(_00638_),
    .A(net3949));
 sg13g2_inv_1 _12084_ (.Y(_00639_),
    .A(net3950));
 sg13g2_inv_1 _12085_ (.Y(_00640_),
    .A(net3950));
 sg13g2_inv_1 _12086_ (.Y(_00641_),
    .A(net3949));
 sg13g2_inv_1 _12087_ (.Y(_00642_),
    .A(net3950));
 sg13g2_inv_1 _12088_ (.Y(_00643_),
    .A(net3951));
 sg13g2_inv_1 _12089_ (.Y(_00644_),
    .A(net3951));
 sg13g2_inv_1 _12090_ (.Y(_00645_),
    .A(net3949));
 sg13g2_inv_1 _12091_ (.Y(_00646_),
    .A(net3947));
 sg13g2_inv_1 _12092_ (.Y(_00647_),
    .A(net3947));
 sg13g2_inv_1 _12093_ (.Y(_00648_),
    .A(net3944));
 sg13g2_inv_1 _12094_ (.Y(_00649_),
    .A(net3946));
 sg13g2_inv_1 _12095_ (.Y(_00650_),
    .A(net3945));
 sg13g2_inv_1 _12096_ (.Y(_00651_),
    .A(net3943));
 sg13g2_inv_1 _12097_ (.Y(_00652_),
    .A(net3943));
 sg13g2_inv_1 _12098_ (.Y(_00653_),
    .A(net3944));
 sg13g2_inv_1 _12099_ (.Y(_00654_),
    .A(net3951));
 sg13g2_inv_1 _12100_ (.Y(_00655_),
    .A(net3946));
 sg13g2_inv_1 _12101_ (.Y(_00656_),
    .A(net3948));
 sg13g2_inv_1 _12102_ (.Y(_00657_),
    .A(net3945));
 sg13g2_inv_1 _12103_ (.Y(_00658_),
    .A(net3943));
 sg13g2_inv_1 _12104_ (.Y(_00659_),
    .A(net3943));
 sg13g2_inv_1 _12105_ (.Y(_00660_),
    .A(net3942));
 sg13g2_inv_1 _12106_ (.Y(_00661_),
    .A(net3942));
 sg13g2_inv_1 _12107_ (.Y(_00662_),
    .A(net3940));
 sg13g2_inv_1 _12108_ (.Y(_00663_),
    .A(net3944));
 sg13g2_inv_1 _12109_ (.Y(_00664_),
    .A(net3947));
 sg13g2_inv_1 _12110_ (.Y(_00665_),
    .A(net3946));
 sg13g2_inv_1 _12111_ (.Y(_00666_),
    .A(net3946));
 sg13g2_inv_1 _12112_ (.Y(_00667_),
    .A(net3946));
 sg13g2_inv_1 _12113_ (.Y(_00668_),
    .A(net3949));
 sg13g2_inv_1 _12114_ (.Y(_00669_),
    .A(net3950));
 sg13g2_inv_1 _12115_ (.Y(_00670_),
    .A(net3949));
 sg13g2_inv_1 _12116_ (.Y(_00671_),
    .A(net3949));
 sg13g2_inv_1 _12117_ (.Y(_00672_),
    .A(net3950));
 sg13g2_inv_1 _12118_ (.Y(_00673_),
    .A(net3951));
 sg13g2_inv_1 _12119_ (.Y(_00674_),
    .A(net3951));
 sg13g2_inv_1 _12120_ (.Y(_00675_),
    .A(net3949));
 sg13g2_inv_1 _12121_ (.Y(_00676_),
    .A(net3947));
 sg13g2_inv_1 _12122_ (.Y(_00677_),
    .A(net3947));
 sg13g2_inv_1 _12123_ (.Y(_00678_),
    .A(net3944));
 sg13g2_inv_1 _12124_ (.Y(_00679_),
    .A(net3946));
 sg13g2_inv_1 _12125_ (.Y(_00680_),
    .A(net3944));
 sg13g2_inv_1 _12126_ (.Y(_00681_),
    .A(net3943));
 sg13g2_inv_1 _12127_ (.Y(_00682_),
    .A(net3943));
 sg13g2_inv_1 _12128_ (.Y(_00683_),
    .A(net3944));
 sg13g2_inv_1 _12129_ (.Y(_00684_),
    .A(net3947));
 sg13g2_inv_1 _12130_ (.Y(_00685_),
    .A(net3948));
 sg13g2_inv_1 _12131_ (.Y(_00686_),
    .A(net3947));
 sg13g2_inv_1 _12132_ (.Y(_00687_),
    .A(net3943));
 sg13g2_inv_1 _12133_ (.Y(_00688_),
    .A(net3946));
 sg13g2_inv_1 _12134_ (.Y(_00689_),
    .A(net3943));
 sg13g2_inv_1 _12135_ (.Y(_00690_),
    .A(net3941));
 sg13g2_inv_1 _12136_ (.Y(_00692_),
    .A(net3940));
 sg13g2_inv_1 _12137_ (.Y(_00693_),
    .A(net3940));
 sg13g2_inv_1 _12138_ (.Y(_00694_),
    .A(net3940));
 sg13g2_dfrbp_1 _12139_ (.CLK(net3840),
    .RESET_B(net418),
    .D(_00695_),
    .Q_N(_00541_),
    .Q(\cpu.regs[13][0] ));
 sg13g2_dfrbp_1 _12140_ (.CLK(net3841),
    .RESET_B(net327),
    .D(_00696_),
    .Q_N(_00540_),
    .Q(\cpu.regs[13][1] ));
 sg13g2_dfrbp_1 _12141_ (.CLK(net3793),
    .RESET_B(net326),
    .D(_00697_),
    .Q_N(_00539_),
    .Q(\cpu.regs[13][2] ));
 sg13g2_dfrbp_1 _12142_ (.CLK(net3862),
    .RESET_B(net325),
    .D(_00698_),
    .Q_N(_00538_),
    .Q(\cpu.regs[13][3] ));
 sg13g2_dfrbp_1 _12143_ (.CLK(net3793),
    .RESET_B(net324),
    .D(_00699_),
    .Q_N(_00537_),
    .Q(\cpu.regs[13][4] ));
 sg13g2_dfrbp_1 _12144_ (.CLK(net3864),
    .RESET_B(net323),
    .D(_00700_),
    .Q_N(_00536_),
    .Q(\cpu.regs[13][5] ));
 sg13g2_dfrbp_1 _12145_ (.CLK(net3847),
    .RESET_B(net322),
    .D(_00701_),
    .Q_N(_00535_),
    .Q(\cpu.regs[13][6] ));
 sg13g2_dfrbp_1 _12146_ (.CLK(net3861),
    .RESET_B(net321),
    .D(_00702_),
    .Q_N(_00534_),
    .Q(\cpu.regs[13][7] ));
 sg13g2_dfrbp_1 _12147_ (.CLK(net3867),
    .RESET_B(net320),
    .D(_00703_),
    .Q_N(_00533_),
    .Q(\cpu.regs[13][8] ));
 sg13g2_dfrbp_1 _12148_ (.CLK(net3854),
    .RESET_B(net319),
    .D(_00704_),
    .Q_N(_00532_),
    .Q(\cpu.regs[13][9] ));
 sg13g2_dfrbp_1 _12149_ (.CLK(net3858),
    .RESET_B(net318),
    .D(_00705_),
    .Q_N(_00531_),
    .Q(\cpu.regs[13][10] ));
 sg13g2_dfrbp_1 _12150_ (.CLK(net3857),
    .RESET_B(net317),
    .D(_00706_),
    .Q_N(_00530_),
    .Q(\cpu.regs[13][11] ));
 sg13g2_dfrbp_1 _12151_ (.CLK(net3804),
    .RESET_B(net316),
    .D(_00707_),
    .Q_N(_00529_),
    .Q(\cpu.regs[13][12] ));
 sg13g2_dfrbp_1 _12152_ (.CLK(net3807),
    .RESET_B(net315),
    .D(_00708_),
    .Q_N(_00528_),
    .Q(\cpu.regs[13][13] ));
 sg13g2_dfrbp_1 _12153_ (.CLK(net3836),
    .RESET_B(net314),
    .D(_00709_),
    .Q_N(_00527_),
    .Q(\cpu.regs[13][14] ));
 sg13g2_dfrbp_1 _12154_ (.CLK(net3851),
    .RESET_B(net313),
    .D(_00710_),
    .Q_N(_00526_),
    .Q(\cpu.regs[13][15] ));
 sg13g2_dfrbp_1 _12155_ (.CLK(net3837),
    .RESET_B(net312),
    .D(_00711_),
    .Q_N(_00525_),
    .Q(\cpu.regs[13][16] ));
 sg13g2_dfrbp_1 _12156_ (.CLK(net3858),
    .RESET_B(net311),
    .D(_00712_),
    .Q_N(_00524_),
    .Q(\cpu.regs[13][17] ));
 sg13g2_dfrbp_1 _12157_ (.CLK(net3830),
    .RESET_B(net310),
    .D(_00713_),
    .Q_N(_00523_),
    .Q(\cpu.regs[13][18] ));
 sg13g2_dfrbp_1 _12158_ (.CLK(net3860),
    .RESET_B(net309),
    .D(_00714_),
    .Q_N(_00522_),
    .Q(\cpu.regs[13][19] ));
 sg13g2_dfrbp_1 _12159_ (.CLK(net3805),
    .RESET_B(net308),
    .D(_00715_),
    .Q_N(_00521_),
    .Q(\cpu.regs[13][20] ));
 sg13g2_dfrbp_1 _12160_ (.CLK(net3822),
    .RESET_B(net307),
    .D(_00716_),
    .Q_N(_00520_),
    .Q(\cpu.regs[13][21] ));
 sg13g2_dfrbp_1 _12161_ (.CLK(net3814),
    .RESET_B(net306),
    .D(_00717_),
    .Q_N(_00519_),
    .Q(\cpu.regs[13][22] ));
 sg13g2_dfrbp_1 _12162_ (.CLK(net3814),
    .RESET_B(net305),
    .D(_00718_),
    .Q_N(_00518_),
    .Q(\cpu.regs[13][23] ));
 sg13g2_dfrbp_1 _12163_ (.CLK(net3816),
    .RESET_B(net304),
    .D(_00719_),
    .Q_N(_00517_),
    .Q(\cpu.regs[13][24] ));
 sg13g2_dfrbp_1 _12164_ (.CLK(net3829),
    .RESET_B(net303),
    .D(_00720_),
    .Q_N(_00516_),
    .Q(\cpu.regs[13][25] ));
 sg13g2_dfrbp_1 _12165_ (.CLK(net3805),
    .RESET_B(net302),
    .D(_00721_),
    .Q_N(_00515_),
    .Q(\cpu.regs[13][26] ));
 sg13g2_dfrbp_1 _12166_ (.CLK(net3825),
    .RESET_B(net301),
    .D(_00722_),
    .Q_N(_00514_),
    .Q(\cpu.regs[13][27] ));
 sg13g2_dfrbp_1 _12167_ (.CLK(net3816),
    .RESET_B(net300),
    .D(_00723_),
    .Q_N(_00513_),
    .Q(\cpu.regs[13][28] ));
 sg13g2_dfrbp_1 _12168_ (.CLK(net3827),
    .RESET_B(net299),
    .D(_00724_),
    .Q_N(_00512_),
    .Q(\cpu.regs[13][29] ));
 sg13g2_dfrbp_1 _12169_ (.CLK(net3809),
    .RESET_B(net298),
    .D(_00725_),
    .Q_N(_00511_),
    .Q(\cpu.regs[13][30] ));
 sg13g2_dfrbp_1 _12170_ (.CLK(net3815),
    .RESET_B(net297),
    .D(_00726_),
    .Q_N(_00510_),
    .Q(\cpu.regs[13][31] ));
 sg13g2_dfrbp_1 _12171_ (.CLK(net3753),
    .RESET_B(net296),
    .D(_00727_),
    .Q_N(_06028_),
    .Q(\irqvect[1][0] ));
 sg13g2_dfrbp_1 _12172_ (.CLK(net3753),
    .RESET_B(net295),
    .D(_00728_),
    .Q_N(_06027_),
    .Q(\irqvect[1][1] ));
 sg13g2_dfrbp_1 _12173_ (.CLK(net3752),
    .RESET_B(net294),
    .D(_00729_),
    .Q_N(_06026_),
    .Q(\irqvect[1][2] ));
 sg13g2_dfrbp_1 _12174_ (.CLK(net3779),
    .RESET_B(net293),
    .D(_00730_),
    .Q_N(_06025_),
    .Q(\irqvect[1][3] ));
 sg13g2_dfrbp_1 _12175_ (.CLK(net3779),
    .RESET_B(net292),
    .D(_00731_),
    .Q_N(_06024_),
    .Q(\irqvect[1][4] ));
 sg13g2_dfrbp_1 _12176_ (.CLK(net3753),
    .RESET_B(net291),
    .D(_00732_),
    .Q_N(_06023_),
    .Q(\irqvect[1][5] ));
 sg13g2_dfrbp_1 _12177_ (.CLK(net3780),
    .RESET_B(net290),
    .D(_00733_),
    .Q_N(_06022_),
    .Q(\irqvect[1][6] ));
 sg13g2_dfrbp_1 _12178_ (.CLK(net3754),
    .RESET_B(net289),
    .D(_00734_),
    .Q_N(_06021_),
    .Q(\irqvect[1][7] ));
 sg13g2_dfrbp_1 _12179_ (.CLK(net3760),
    .RESET_B(net288),
    .D(_00735_),
    .Q_N(_06020_),
    .Q(\irqvect[1][8] ));
 sg13g2_dfrbp_1 _12180_ (.CLK(net3746),
    .RESET_B(net287),
    .D(_00736_),
    .Q_N(_06019_),
    .Q(\irqvect[1][9] ));
 sg13g2_dfrbp_1 _12181_ (.CLK(net3756),
    .RESET_B(net286),
    .D(_00737_),
    .Q_N(_06018_),
    .Q(\irqvect[1][10] ));
 sg13g2_dfrbp_1 _12182_ (.CLK(net3742),
    .RESET_B(net285),
    .D(_00738_),
    .Q_N(_06017_),
    .Q(\irqvect[1][11] ));
 sg13g2_dfrbp_1 _12183_ (.CLK(net3745),
    .RESET_B(net284),
    .D(_00739_),
    .Q_N(_06016_),
    .Q(\irqvect[1][12] ));
 sg13g2_dfrbp_1 _12184_ (.CLK(net3758),
    .RESET_B(net283),
    .D(_00740_),
    .Q_N(_06015_),
    .Q(\irqvect[1][13] ));
 sg13g2_dfrbp_1 _12185_ (.CLK(net3750),
    .RESET_B(net282),
    .D(_00741_),
    .Q_N(_06014_),
    .Q(\irqvect[1][14] ));
 sg13g2_dfrbp_1 _12186_ (.CLK(net3751),
    .RESET_B(net281),
    .D(_00742_),
    .Q_N(_06013_),
    .Q(\irqvect[1][15] ));
 sg13g2_dfrbp_1 _12187_ (.CLK(net3750),
    .RESET_B(net280),
    .D(_00743_),
    .Q_N(_06012_),
    .Q(\irqvect[1][16] ));
 sg13g2_dfrbp_1 _12188_ (.CLK(net3745),
    .RESET_B(net279),
    .D(_00744_),
    .Q_N(_06011_),
    .Q(\irqvect[1][17] ));
 sg13g2_dfrbp_1 _12189_ (.CLK(net3744),
    .RESET_B(net278),
    .D(_00745_),
    .Q_N(_06010_),
    .Q(\irqvect[1][18] ));
 sg13g2_dfrbp_1 _12190_ (.CLK(net3749),
    .RESET_B(net277),
    .D(_00746_),
    .Q_N(_06009_),
    .Q(\irqvect[1][19] ));
 sg13g2_dfrbp_1 _12191_ (.CLK(net3745),
    .RESET_B(net276),
    .D(_00747_),
    .Q_N(_06008_),
    .Q(\irqvect[1][20] ));
 sg13g2_dfrbp_1 _12192_ (.CLK(net3746),
    .RESET_B(net275),
    .D(_00748_),
    .Q_N(_06007_),
    .Q(\irqvect[1][21] ));
 sg13g2_dfrbp_1 _12193_ (.CLK(net3743),
    .RESET_B(net274),
    .D(_00749_),
    .Q_N(_06006_),
    .Q(\irqvect[1][22] ));
 sg13g2_dfrbp_1 _12194_ (.CLK(net3762),
    .RESET_B(net273),
    .D(_00750_),
    .Q_N(_06005_),
    .Q(\irqvect[1][23] ));
 sg13g2_dfrbp_1 _12195_ (.CLK(net3743),
    .RESET_B(net272),
    .D(_00751_),
    .Q_N(_06004_),
    .Q(\irqvect[1][24] ));
 sg13g2_dfrbp_1 _12196_ (.CLK(net3756),
    .RESET_B(net271),
    .D(_00752_),
    .Q_N(_06003_),
    .Q(\irqvect[1][25] ));
 sg13g2_dfrbp_1 _12197_ (.CLK(net3744),
    .RESET_B(net270),
    .D(_00753_),
    .Q_N(_06002_),
    .Q(\irqvect[1][26] ));
 sg13g2_dfrbp_1 _12198_ (.CLK(net3747),
    .RESET_B(net269),
    .D(_00754_),
    .Q_N(_06001_),
    .Q(\irqvect[1][27] ));
 sg13g2_dfrbp_1 _12199_ (.CLK(net3740),
    .RESET_B(net268),
    .D(_00755_),
    .Q_N(_06000_),
    .Q(\irqvect[1][28] ));
 sg13g2_dfrbp_1 _12200_ (.CLK(net3740),
    .RESET_B(net267),
    .D(_00756_),
    .Q_N(_05999_),
    .Q(\irqvect[1][29] ));
 sg13g2_dfrbp_1 _12201_ (.CLK(net3792),
    .RESET_B(net266),
    .D(_00757_),
    .Q_N(_00509_),
    .Q(\cpu.regs[1][0] ));
 sg13g2_dfrbp_1 _12202_ (.CLK(net3843),
    .RESET_B(net265),
    .D(_00758_),
    .Q_N(_00508_),
    .Q(\cpu.regs[1][1] ));
 sg13g2_dfrbp_1 _12203_ (.CLK(net3796),
    .RESET_B(net264),
    .D(_00759_),
    .Q_N(_00507_),
    .Q(\cpu.regs[1][2] ));
 sg13g2_dfrbp_1 _12204_ (.CLK(net3849),
    .RESET_B(net263),
    .D(_00760_),
    .Q_N(_00506_),
    .Q(\cpu.regs[1][3] ));
 sg13g2_dfrbp_1 _12205_ (.CLK(net3794),
    .RESET_B(net262),
    .D(_00761_),
    .Q_N(_00505_),
    .Q(\cpu.regs[1][4] ));
 sg13g2_dfrbp_1 _12206_ (.CLK(net3863),
    .RESET_B(net261),
    .D(_00762_),
    .Q_N(_00504_),
    .Q(\cpu.regs[1][5] ));
 sg13g2_dfrbp_1 _12207_ (.CLK(net3843),
    .RESET_B(net260),
    .D(_00763_),
    .Q_N(_00503_),
    .Q(\cpu.regs[1][6] ));
 sg13g2_dfrbp_1 _12208_ (.CLK(net3848),
    .RESET_B(net259),
    .D(_00764_),
    .Q_N(_00502_),
    .Q(\cpu.regs[1][7] ));
 sg13g2_dfrbp_1 _12209_ (.CLK(net3863),
    .RESET_B(net258),
    .D(_00765_),
    .Q_N(_00501_),
    .Q(\cpu.regs[1][8] ));
 sg13g2_dfrbp_1 _12210_ (.CLK(net3836),
    .RESET_B(net257),
    .D(_00766_),
    .Q_N(_00500_),
    .Q(\cpu.regs[1][9] ));
 sg13g2_dfrbp_1 _12211_ (.CLK(net3867),
    .RESET_B(net256),
    .D(_00767_),
    .Q_N(_00499_),
    .Q(\cpu.regs[1][10] ));
 sg13g2_dfrbp_1 _12212_ (.CLK(net3856),
    .RESET_B(net255),
    .D(_00768_),
    .Q_N(_00498_),
    .Q(\cpu.regs[1][11] ));
 sg13g2_dfrbp_1 _12213_ (.CLK(net3799),
    .RESET_B(net254),
    .D(_00769_),
    .Q_N(_00497_),
    .Q(\cpu.regs[1][12] ));
 sg13g2_dfrbp_1 _12214_ (.CLK(net3768),
    .RESET_B(net253),
    .D(_00770_),
    .Q_N(_00496_),
    .Q(\cpu.regs[1][13] ));
 sg13g2_dfrbp_1 _12215_ (.CLK(net3851),
    .RESET_B(net252),
    .D(_00771_),
    .Q_N(_00495_),
    .Q(\cpu.regs[1][14] ));
 sg13g2_dfrbp_1 _12216_ (.CLK(net3834),
    .RESET_B(net251),
    .D(_00772_),
    .Q_N(_00494_),
    .Q(\cpu.regs[1][15] ));
 sg13g2_dfrbp_1 _12217_ (.CLK(net3846),
    .RESET_B(net250),
    .D(_00773_),
    .Q_N(_00493_),
    .Q(\cpu.regs[1][16] ));
 sg13g2_dfrbp_1 _12218_ (.CLK(net3858),
    .RESET_B(net249),
    .D(_00774_),
    .Q_N(_00492_),
    .Q(\cpu.regs[1][17] ));
 sg13g2_dfrbp_1 _12219_ (.CLK(net3828),
    .RESET_B(net248),
    .D(_00775_),
    .Q_N(_00491_),
    .Q(\cpu.regs[1][18] ));
 sg13g2_dfrbp_1 _12220_ (.CLK(net3856),
    .RESET_B(net247),
    .D(_00776_),
    .Q_N(_00490_),
    .Q(\cpu.regs[1][19] ));
 sg13g2_dfrbp_1 _12221_ (.CLK(net3800),
    .RESET_B(net246),
    .D(_00777_),
    .Q_N(_00489_),
    .Q(\cpu.regs[1][20] ));
 sg13g2_dfrbp_1 _12222_ (.CLK(net3819),
    .RESET_B(net245),
    .D(_00778_),
    .Q_N(_00488_),
    .Q(\cpu.regs[1][21] ));
 sg13g2_dfrbp_1 _12223_ (.CLK(net3820),
    .RESET_B(net244),
    .D(_00779_),
    .Q_N(_00487_),
    .Q(\cpu.regs[1][22] ));
 sg13g2_dfrbp_1 _12224_ (.CLK(net3820),
    .RESET_B(net243),
    .D(_00780_),
    .Q_N(_00486_),
    .Q(\cpu.regs[1][23] ));
 sg13g2_dfrbp_1 _12225_ (.CLK(net3810),
    .RESET_B(net242),
    .D(_00781_),
    .Q_N(_00485_),
    .Q(\cpu.regs[1][24] ));
 sg13g2_dfrbp_1 _12226_ (.CLK(net3828),
    .RESET_B(net241),
    .D(_00782_),
    .Q_N(_00484_),
    .Q(\cpu.regs[1][25] ));
 sg13g2_dfrbp_1 _12227_ (.CLK(net3800),
    .RESET_B(net240),
    .D(_00783_),
    .Q_N(_00483_),
    .Q(\cpu.regs[1][26] ));
 sg13g2_dfrbp_1 _12228_ (.CLK(net3825),
    .RESET_B(net239),
    .D(_00784_),
    .Q_N(_00482_),
    .Q(\cpu.regs[1][27] ));
 sg13g2_dfrbp_1 _12229_ (.CLK(net3812),
    .RESET_B(net238),
    .D(_00785_),
    .Q_N(_00481_),
    .Q(\cpu.regs[1][28] ));
 sg13g2_dfrbp_1 _12230_ (.CLK(net3827),
    .RESET_B(net237),
    .D(_00786_),
    .Q_N(_00480_),
    .Q(\cpu.regs[1][29] ));
 sg13g2_dfrbp_1 _12231_ (.CLK(net3767),
    .RESET_B(net236),
    .D(_00787_),
    .Q_N(_00479_),
    .Q(\cpu.regs[1][30] ));
 sg13g2_dfrbp_1 _12232_ (.CLK(net3799),
    .RESET_B(net235),
    .D(_00788_),
    .Q_N(_00478_),
    .Q(\cpu.regs[1][31] ));
 sg13g2_dfrbp_1 _12233_ (.CLK(net3840),
    .RESET_B(net234),
    .D(_00789_),
    .Q_N(_00477_),
    .Q(\cpu.regs[11][0] ));
 sg13g2_dfrbp_1 _12234_ (.CLK(net3843),
    .RESET_B(net233),
    .D(_00790_),
    .Q_N(_00476_),
    .Q(\cpu.regs[11][1] ));
 sg13g2_dfrbp_1 _12235_ (.CLK(net3795),
    .RESET_B(net232),
    .D(_00791_),
    .Q_N(_00475_),
    .Q(\cpu.regs[11][2] ));
 sg13g2_dfrbp_1 _12236_ (.CLK(net3862),
    .RESET_B(net231),
    .D(_00792_),
    .Q_N(_00474_),
    .Q(\cpu.regs[11][3] ));
 sg13g2_dfrbp_1 _12237_ (.CLK(net3844),
    .RESET_B(net230),
    .D(_00793_),
    .Q_N(_00473_),
    .Q(\cpu.regs[11][4] ));
 sg13g2_dfrbp_1 _12238_ (.CLK(net3864),
    .RESET_B(net229),
    .D(_00794_),
    .Q_N(_00472_),
    .Q(\cpu.regs[11][5] ));
 sg13g2_dfrbp_1 _12239_ (.CLK(net3847),
    .RESET_B(net228),
    .D(_00795_),
    .Q_N(_00471_),
    .Q(\cpu.regs[11][6] ));
 sg13g2_dfrbp_1 _12240_ (.CLK(net3864),
    .RESET_B(net227),
    .D(_00796_),
    .Q_N(_00470_),
    .Q(\cpu.regs[11][7] ));
 sg13g2_dfrbp_1 _12241_ (.CLK(net3868),
    .RESET_B(net226),
    .D(_00797_),
    .Q_N(_00469_),
    .Q(\cpu.regs[11][8] ));
 sg13g2_dfrbp_1 _12242_ (.CLK(net3845),
    .RESET_B(net225),
    .D(_00798_),
    .Q_N(_00468_),
    .Q(\cpu.regs[11][9] ));
 sg13g2_dfrbp_1 _12243_ (.CLK(net3859),
    .RESET_B(net224),
    .D(_00799_),
    .Q_N(_00467_),
    .Q(\cpu.regs[11][10] ));
 sg13g2_dfrbp_1 _12244_ (.CLK(net3857),
    .RESET_B(net223),
    .D(_00800_),
    .Q_N(_00466_),
    .Q(\cpu.regs[11][11] ));
 sg13g2_dfrbp_1 _12245_ (.CLK(net3807),
    .RESET_B(net222),
    .D(_00801_),
    .Q_N(_00465_),
    .Q(\cpu.regs[11][12] ));
 sg13g2_dfrbp_1 _12246_ (.CLK(net3808),
    .RESET_B(net221),
    .D(_00802_),
    .Q_N(_00464_),
    .Q(\cpu.regs[11][13] ));
 sg13g2_dfrbp_1 _12247_ (.CLK(net3854),
    .RESET_B(net220),
    .D(_00803_),
    .Q_N(_00463_),
    .Q(\cpu.regs[11][14] ));
 sg13g2_dfrbp_1 _12248_ (.CLK(net3852),
    .RESET_B(net219),
    .D(_00804_),
    .Q_N(_00462_),
    .Q(\cpu.regs[11][15] ));
 sg13g2_dfrbp_1 _12249_ (.CLK(net3837),
    .RESET_B(net218),
    .D(_00805_),
    .Q_N(_00461_),
    .Q(\cpu.regs[11][16] ));
 sg13g2_dfrbp_1 _12250_ (.CLK(net3859),
    .RESET_B(net217),
    .D(_00806_),
    .Q_N(_00460_),
    .Q(\cpu.regs[11][17] ));
 sg13g2_dfrbp_1 _12251_ (.CLK(net3860),
    .RESET_B(net216),
    .D(_00807_),
    .Q_N(_00459_),
    .Q(\cpu.regs[11][18] ));
 sg13g2_dfrbp_1 _12252_ (.CLK(net3830),
    .RESET_B(net215),
    .D(_00808_),
    .Q_N(_00458_),
    .Q(\cpu.regs[11][19] ));
 sg13g2_dfrbp_1 _12253_ (.CLK(net3803),
    .RESET_B(net214),
    .D(_00809_),
    .Q_N(_00457_),
    .Q(\cpu.regs[11][20] ));
 sg13g2_dfrbp_1 _12254_ (.CLK(net3819),
    .RESET_B(net213),
    .D(_00810_),
    .Q_N(_00456_),
    .Q(\cpu.regs[11][21] ));
 sg13g2_dfrbp_1 _12255_ (.CLK(net3814),
    .RESET_B(net212),
    .D(_00811_),
    .Q_N(_00455_),
    .Q(\cpu.regs[11][22] ));
 sg13g2_dfrbp_1 _12256_ (.CLK(net3818),
    .RESET_B(net211),
    .D(_00812_),
    .Q_N(_00454_),
    .Q(\cpu.regs[11][23] ));
 sg13g2_dfrbp_1 _12257_ (.CLK(net3813),
    .RESET_B(net210),
    .D(_00813_),
    .Q_N(_00453_),
    .Q(\cpu.regs[11][24] ));
 sg13g2_dfrbp_1 _12258_ (.CLK(net3829),
    .RESET_B(net209),
    .D(_00814_),
    .Q_N(_00452_),
    .Q(\cpu.regs[11][25] ));
 sg13g2_dfrbp_1 _12259_ (.CLK(net3804),
    .RESET_B(net208),
    .D(_00815_),
    .Q_N(_00451_),
    .Q(\cpu.regs[11][26] ));
 sg13g2_dfrbp_1 _12260_ (.CLK(net3817),
    .RESET_B(net207),
    .D(_00816_),
    .Q_N(_00450_),
    .Q(\cpu.regs[11][27] ));
 sg13g2_dfrbp_1 _12261_ (.CLK(net3816),
    .RESET_B(net206),
    .D(_00817_),
    .Q_N(_00449_),
    .Q(\cpu.regs[11][28] ));
 sg13g2_dfrbp_1 _12262_ (.CLK(net3826),
    .RESET_B(net205),
    .D(_00818_),
    .Q_N(_00448_),
    .Q(\cpu.regs[11][29] ));
 sg13g2_dfrbp_1 _12263_ (.CLK(net3809),
    .RESET_B(net204),
    .D(_00819_),
    .Q_N(_00447_),
    .Q(\cpu.regs[11][30] ));
 sg13g2_dfrbp_1 _12264_ (.CLK(net3802),
    .RESET_B(net203),
    .D(_00820_),
    .Q_N(_00446_),
    .Q(\cpu.regs[11][31] ));
 sg13g2_dfrbp_1 _12265_ (.CLK(net3840),
    .RESET_B(net202),
    .D(_00821_),
    .Q_N(_00445_),
    .Q(\cpu.regs[12][0] ));
 sg13g2_dfrbp_1 _12266_ (.CLK(net3841),
    .RESET_B(net201),
    .D(_00822_),
    .Q_N(_00444_),
    .Q(\cpu.regs[12][1] ));
 sg13g2_dfrbp_1 _12267_ (.CLK(net3795),
    .RESET_B(net200),
    .D(_00823_),
    .Q_N(_00443_),
    .Q(\cpu.regs[12][2] ));
 sg13g2_dfrbp_1 _12268_ (.CLK(net3861),
    .RESET_B(net199),
    .D(_00824_),
    .Q_N(_00442_),
    .Q(\cpu.regs[12][3] ));
 sg13g2_dfrbp_1 _12269_ (.CLK(net3793),
    .RESET_B(net198),
    .D(_00825_),
    .Q_N(_00441_),
    .Q(\cpu.regs[12][4] ));
 sg13g2_dfrbp_1 _12270_ (.CLK(net3864),
    .RESET_B(net197),
    .D(_00826_),
    .Q_N(_00440_),
    .Q(\cpu.regs[12][5] ));
 sg13g2_dfrbp_1 _12271_ (.CLK(net3847),
    .RESET_B(net196),
    .D(_00827_),
    .Q_N(_00439_),
    .Q(\cpu.regs[12][6] ));
 sg13g2_dfrbp_1 _12272_ (.CLK(net3864),
    .RESET_B(net195),
    .D(_00828_),
    .Q_N(_00438_),
    .Q(\cpu.regs[12][7] ));
 sg13g2_dfrbp_1 _12273_ (.CLK(net3867),
    .RESET_B(net194),
    .D(_00829_),
    .Q_N(_00437_),
    .Q(\cpu.regs[12][8] ));
 sg13g2_dfrbp_1 _12274_ (.CLK(net3836),
    .RESET_B(net193),
    .D(_00830_),
    .Q_N(_00436_),
    .Q(\cpu.regs[12][9] ));
 sg13g2_dfrbp_1 _12275_ (.CLK(net3867),
    .RESET_B(net192),
    .D(_00831_),
    .Q_N(_00435_),
    .Q(\cpu.regs[12][10] ));
 sg13g2_dfrbp_1 _12276_ (.CLK(net3857),
    .RESET_B(net191),
    .D(_00832_),
    .Q_N(_00434_),
    .Q(\cpu.regs[12][11] ));
 sg13g2_dfrbp_1 _12277_ (.CLK(net3804),
    .RESET_B(net190),
    .D(_00833_),
    .Q_N(_00433_),
    .Q(\cpu.regs[12][12] ));
 sg13g2_dfrbp_1 _12278_ (.CLK(net3805),
    .RESET_B(net189),
    .D(_00834_),
    .Q_N(_00432_),
    .Q(\cpu.regs[12][13] ));
 sg13g2_dfrbp_1 _12279_ (.CLK(net3836),
    .RESET_B(net188),
    .D(_00835_),
    .Q_N(_00431_),
    .Q(\cpu.regs[12][14] ));
 sg13g2_dfrbp_1 _12280_ (.CLK(net3851),
    .RESET_B(net187),
    .D(_00836_),
    .Q_N(_00430_),
    .Q(\cpu.regs[12][15] ));
 sg13g2_dfrbp_1 _12281_ (.CLK(net3837),
    .RESET_B(net186),
    .D(_00837_),
    .Q_N(_00429_),
    .Q(\cpu.regs[12][16] ));
 sg13g2_dfrbp_1 _12282_ (.CLK(net3858),
    .RESET_B(net185),
    .D(_00838_),
    .Q_N(_00428_),
    .Q(\cpu.regs[12][17] ));
 sg13g2_dfrbp_1 _12283_ (.CLK(net3830),
    .RESET_B(net184),
    .D(_00839_),
    .Q_N(_00427_),
    .Q(\cpu.regs[12][18] ));
 sg13g2_dfrbp_1 _12284_ (.CLK(net3831),
    .RESET_B(net183),
    .D(_00840_),
    .Q_N(_00426_),
    .Q(\cpu.regs[12][19] ));
 sg13g2_dfrbp_1 _12285_ (.CLK(net3803),
    .RESET_B(net182),
    .D(_00841_),
    .Q_N(_00425_),
    .Q(\cpu.regs[12][20] ));
 sg13g2_dfrbp_1 _12286_ (.CLK(net3819),
    .RESET_B(net181),
    .D(_00842_),
    .Q_N(_00424_),
    .Q(\cpu.regs[12][21] ));
 sg13g2_dfrbp_1 _12287_ (.CLK(net3815),
    .RESET_B(net180),
    .D(_00843_),
    .Q_N(_00423_),
    .Q(\cpu.regs[12][22] ));
 sg13g2_dfrbp_1 _12288_ (.CLK(net3818),
    .RESET_B(net179),
    .D(_00844_),
    .Q_N(_00422_),
    .Q(\cpu.regs[12][23] ));
 sg13g2_dfrbp_1 _12289_ (.CLK(net3816),
    .RESET_B(net178),
    .D(_00845_),
    .Q_N(_00421_),
    .Q(\cpu.regs[12][24] ));
 sg13g2_dfrbp_1 _12290_ (.CLK(net3821),
    .RESET_B(net177),
    .D(_00846_),
    .Q_N(_00420_),
    .Q(\cpu.regs[12][25] ));
 sg13g2_dfrbp_1 _12291_ (.CLK(net3803),
    .RESET_B(net176),
    .D(_00847_),
    .Q_N(_00419_),
    .Q(\cpu.regs[12][26] ));
 sg13g2_dfrbp_1 _12292_ (.CLK(net3817),
    .RESET_B(net175),
    .D(_00848_),
    .Q_N(_00418_),
    .Q(\cpu.regs[12][27] ));
 sg13g2_dfrbp_1 _12293_ (.CLK(net3816),
    .RESET_B(net174),
    .D(_00849_),
    .Q_N(_00417_),
    .Q(\cpu.regs[12][28] ));
 sg13g2_dfrbp_1 _12294_ (.CLK(net3827),
    .RESET_B(net173),
    .D(_00850_),
    .Q_N(_00416_),
    .Q(\cpu.regs[12][29] ));
 sg13g2_dfrbp_1 _12295_ (.CLK(net3809),
    .RESET_B(net172),
    .D(_00851_),
    .Q_N(_00415_),
    .Q(\cpu.regs[12][30] ));
 sg13g2_dfrbp_1 _12296_ (.CLK(net3815),
    .RESET_B(net171),
    .D(_00852_),
    .Q_N(_00414_),
    .Q(\cpu.regs[12][31] ));
 sg13g2_dfrbp_1 _12297_ (.CLK(net3794),
    .RESET_B(net170),
    .D(_00853_),
    .Q_N(_00413_),
    .Q(\cpu.regs[7][0] ));
 sg13g2_dfrbp_1 _12298_ (.CLK(net3842),
    .RESET_B(net169),
    .D(_00854_),
    .Q_N(_00412_),
    .Q(\cpu.regs[7][1] ));
 sg13g2_dfrbp_1 _12299_ (.CLK(net3793),
    .RESET_B(net168),
    .D(_00855_),
    .Q_N(_00411_),
    .Q(\cpu.regs[7][2] ));
 sg13g2_dfrbp_1 _12300_ (.CLK(net3846),
    .RESET_B(net167),
    .D(_00856_),
    .Q_N(_00410_),
    .Q(\cpu.regs[7][3] ));
 sg13g2_dfrbp_1 _12301_ (.CLK(net3795),
    .RESET_B(net166),
    .D(_00857_),
    .Q_N(_00409_),
    .Q(\cpu.regs[7][4] ));
 sg13g2_dfrbp_1 _12302_ (.CLK(net3865),
    .RESET_B(net165),
    .D(_00858_),
    .Q_N(_00408_),
    .Q(\cpu.regs[7][5] ));
 sg13g2_dfrbp_1 _12303_ (.CLK(net3843),
    .RESET_B(net164),
    .D(_00859_),
    .Q_N(_00407_),
    .Q(\cpu.regs[7][6] ));
 sg13g2_dfrbp_1 _12304_ (.CLK(net3848),
    .RESET_B(net163),
    .D(_00860_),
    .Q_N(_00406_),
    .Q(\cpu.regs[7][7] ));
 sg13g2_dfrbp_1 _12305_ (.CLK(net3845),
    .RESET_B(net162),
    .D(_00861_),
    .Q_N(_00405_),
    .Q(\cpu.regs[7][8] ));
 sg13g2_dfrbp_1 _12306_ (.CLK(net3834),
    .RESET_B(net161),
    .D(_00862_),
    .Q_N(_00404_),
    .Q(\cpu.regs[7][9] ));
 sg13g2_dfrbp_1 _12307_ (.CLK(net3853),
    .RESET_B(net160),
    .D(_00863_),
    .Q_N(_00403_),
    .Q(\cpu.regs[7][10] ));
 sg13g2_dfrbp_1 _12308_ (.CLK(net3852),
    .RESET_B(net159),
    .D(_00864_),
    .Q_N(_00402_),
    .Q(\cpu.regs[7][11] ));
 sg13g2_dfrbp_1 _12309_ (.CLK(net3761),
    .RESET_B(net158),
    .D(_00865_),
    .Q_N(_00401_),
    .Q(\cpu.regs[7][12] ));
 sg13g2_dfrbp_1 _12310_ (.CLK(net3762),
    .RESET_B(net157),
    .D(_00866_),
    .Q_N(_00400_),
    .Q(\cpu.regs[7][13] ));
 sg13g2_dfrbp_1 _12311_ (.CLK(net3836),
    .RESET_B(net156),
    .D(_00867_),
    .Q_N(_00399_),
    .Q(\cpu.regs[7][14] ));
 sg13g2_dfrbp_1 _12312_ (.CLK(net3835),
    .RESET_B(net155),
    .D(_00868_),
    .Q_N(_00398_),
    .Q(\cpu.regs[7][15] ));
 sg13g2_dfrbp_1 _12313_ (.CLK(net3839),
    .RESET_B(net154),
    .D(_00869_),
    .Q_N(_00397_),
    .Q(\cpu.regs[7][16] ));
 sg13g2_dfrbp_1 _12314_ (.CLK(net3853),
    .RESET_B(net153),
    .D(_00870_),
    .Q_N(_00396_),
    .Q(\cpu.regs[7][17] ));
 sg13g2_dfrbp_1 _12315_ (.CLK(net3831),
    .RESET_B(net152),
    .D(_00871_),
    .Q_N(_00395_),
    .Q(\cpu.regs[7][18] ));
 sg13g2_dfrbp_1 _12316_ (.CLK(net3826),
    .RESET_B(net151),
    .D(_00872_),
    .Q_N(_00394_),
    .Q(\cpu.regs[7][19] ));
 sg13g2_dfrbp_1 _12317_ (.CLK(net3762),
    .RESET_B(net150),
    .D(_00873_),
    .Q_N(_00393_),
    .Q(\cpu.regs[7][20] ));
 sg13g2_dfrbp_1 _12318_ (.CLK(net3818),
    .RESET_B(net149),
    .D(_00874_),
    .Q_N(_00392_),
    .Q(\cpu.regs[7][21] ));
 sg13g2_dfrbp_1 _12319_ (.CLK(net3825),
    .RESET_B(net148),
    .D(_00875_),
    .Q_N(_00391_),
    .Q(\cpu.regs[7][22] ));
 sg13g2_dfrbp_1 _12320_ (.CLK(net3820),
    .RESET_B(net147),
    .D(_00876_),
    .Q_N(_00390_),
    .Q(\cpu.regs[7][23] ));
 sg13g2_dfrbp_1 _12321_ (.CLK(net3806),
    .RESET_B(net146),
    .D(_00877_),
    .Q_N(_00389_),
    .Q(\cpu.regs[7][24] ));
 sg13g2_dfrbp_1 _12322_ (.CLK(net3821),
    .RESET_B(net145),
    .D(_00878_),
    .Q_N(_00388_),
    .Q(\cpu.regs[7][25] ));
 sg13g2_dfrbp_1 _12323_ (.CLK(net3800),
    .RESET_B(net144),
    .D(_00879_),
    .Q_N(_00387_),
    .Q(\cpu.regs[7][26] ));
 sg13g2_dfrbp_1 _12324_ (.CLK(net3824),
    .RESET_B(net143),
    .D(_00880_),
    .Q_N(_00386_),
    .Q(\cpu.regs[7][27] ));
 sg13g2_dfrbp_1 _12325_ (.CLK(net3810),
    .RESET_B(net142),
    .D(_00881_),
    .Q_N(_00385_),
    .Q(\cpu.regs[7][28] ));
 sg13g2_dfrbp_1 _12326_ (.CLK(net3811),
    .RESET_B(net141),
    .D(_00882_),
    .Q_N(_00384_),
    .Q(\cpu.regs[7][29] ));
 sg13g2_dfrbp_1 _12327_ (.CLK(net3763),
    .RESET_B(net140),
    .D(_00883_),
    .Q_N(_00383_),
    .Q(\cpu.regs[7][30] ));
 sg13g2_dfrbp_1 _12328_ (.CLK(net3767),
    .RESET_B(net139),
    .D(_00884_),
    .Q_N(_00382_),
    .Q(\cpu.regs[7][31] ));
 sg13g2_dfrbp_1 _12329_ (.CLK(net3792),
    .RESET_B(net138),
    .D(_00885_),
    .Q_N(_00381_),
    .Q(\cpu.regs[2][0] ));
 sg13g2_dfrbp_1 _12330_ (.CLK(net3842),
    .RESET_B(net137),
    .D(_00886_),
    .Q_N(_00380_),
    .Q(\cpu.regs[2][1] ));
 sg13g2_dfrbp_1 _12331_ (.CLK(net3792),
    .RESET_B(net136),
    .D(_00887_),
    .Q_N(_00379_),
    .Q(\cpu.regs[2][2] ));
 sg13g2_dfrbp_1 _12332_ (.CLK(net3849),
    .RESET_B(net135),
    .D(_00888_),
    .Q_N(_00378_),
    .Q(\cpu.regs[2][3] ));
 sg13g2_dfrbp_1 _12333_ (.CLK(net3794),
    .RESET_B(net134),
    .D(_00889_),
    .Q_N(_00377_),
    .Q(\cpu.regs[2][4] ));
 sg13g2_dfrbp_1 _12334_ (.CLK(net3863),
    .RESET_B(net133),
    .D(_00890_),
    .Q_N(_00376_),
    .Q(\cpu.regs[2][5] ));
 sg13g2_dfrbp_1 _12335_ (.CLK(net3843),
    .RESET_B(net132),
    .D(_00891_),
    .Q_N(_00375_),
    .Q(\cpu.regs[2][6] ));
 sg13g2_dfrbp_1 _12336_ (.CLK(net3848),
    .RESET_B(net131),
    .D(_00892_),
    .Q_N(_00374_),
    .Q(\cpu.regs[2][7] ));
 sg13g2_dfrbp_1 _12337_ (.CLK(net3863),
    .RESET_B(net130),
    .D(_00893_),
    .Q_N(_00373_),
    .Q(\cpu.regs[2][8] ));
 sg13g2_dfrbp_1 _12338_ (.CLK(net3838),
    .RESET_B(net129),
    .D(_00894_),
    .Q_N(_00372_),
    .Q(\cpu.regs[2][9] ));
 sg13g2_dfrbp_1 _12339_ (.CLK(net3861),
    .RESET_B(net128),
    .D(_00895_),
    .Q_N(_00371_),
    .Q(\cpu.regs[2][10] ));
 sg13g2_dfrbp_1 _12340_ (.CLK(net3857),
    .RESET_B(net127),
    .D(_00896_),
    .Q_N(_00370_),
    .Q(\cpu.regs[2][11] ));
 sg13g2_dfrbp_1 _12341_ (.CLK(net3799),
    .RESET_B(net126),
    .D(_00897_),
    .Q_N(_00369_),
    .Q(\cpu.regs[2][12] ));
 sg13g2_dfrbp_1 _12342_ (.CLK(net3768),
    .RESET_B(net125),
    .D(_00898_),
    .Q_N(_00368_),
    .Q(\cpu.regs[2][13] ));
 sg13g2_dfrbp_1 _12343_ (.CLK(net3851),
    .RESET_B(net124),
    .D(_00899_),
    .Q_N(_00367_),
    .Q(\cpu.regs[2][14] ));
 sg13g2_dfrbp_1 _12344_ (.CLK(net3835),
    .RESET_B(net123),
    .D(_00900_),
    .Q_N(_00366_),
    .Q(\cpu.regs[2][15] ));
 sg13g2_dfrbp_1 _12345_ (.CLK(net3841),
    .RESET_B(net122),
    .D(_00901_),
    .Q_N(_00365_),
    .Q(\cpu.regs[2][16] ));
 sg13g2_dfrbp_1 _12346_ (.CLK(net3853),
    .RESET_B(net121),
    .D(_00902_),
    .Q_N(_00364_),
    .Q(\cpu.regs[2][17] ));
 sg13g2_dfrbp_1 _12347_ (.CLK(net3828),
    .RESET_B(net120),
    .D(_00903_),
    .Q_N(_00363_),
    .Q(\cpu.regs[2][18] ));
 sg13g2_dfrbp_1 _12348_ (.CLK(net3831),
    .RESET_B(net119),
    .D(_00904_),
    .Q_N(_00362_),
    .Q(\cpu.regs[2][19] ));
 sg13g2_dfrbp_1 _12349_ (.CLK(net3801),
    .RESET_B(net118),
    .D(_00905_),
    .Q_N(_00361_),
    .Q(\cpu.regs[2][20] ));
 sg13g2_dfrbp_1 _12350_ (.CLK(net3818),
    .RESET_B(net117),
    .D(_00906_),
    .Q_N(_00360_),
    .Q(\cpu.regs[2][21] ));
 sg13g2_dfrbp_1 _12351_ (.CLK(net3828),
    .RESET_B(net116),
    .D(_00907_),
    .Q_N(_00359_),
    .Q(\cpu.regs[2][22] ));
 sg13g2_dfrbp_1 _12352_ (.CLK(net3820),
    .RESET_B(net115),
    .D(_00908_),
    .Q_N(_00358_),
    .Q(\cpu.regs[2][23] ));
 sg13g2_dfrbp_1 _12353_ (.CLK(net3810),
    .RESET_B(net114),
    .D(_00909_),
    .Q_N(_00357_),
    .Q(\cpu.regs[2][24] ));
 sg13g2_dfrbp_1 _12354_ (.CLK(net3828),
    .RESET_B(net113),
    .D(_00910_),
    .Q_N(_00356_),
    .Q(\cpu.regs[2][25] ));
 sg13g2_dfrbp_1 _12355_ (.CLK(net3800),
    .RESET_B(net112),
    .D(_00911_),
    .Q_N(_00355_),
    .Q(\cpu.regs[2][26] ));
 sg13g2_dfrbp_1 _12356_ (.CLK(net3826),
    .RESET_B(net111),
    .D(_00912_),
    .Q_N(_00354_),
    .Q(\cpu.regs[2][27] ));
 sg13g2_dfrbp_1 _12357_ (.CLK(net3812),
    .RESET_B(net110),
    .D(_00913_),
    .Q_N(_00353_),
    .Q(\cpu.regs[2][28] ));
 sg13g2_dfrbp_1 _12358_ (.CLK(net3827),
    .RESET_B(net109),
    .D(_00914_),
    .Q_N(_00352_),
    .Q(\cpu.regs[2][29] ));
 sg13g2_dfrbp_1 _12359_ (.CLK(net3767),
    .RESET_B(net108),
    .D(_00915_),
    .Q_N(_00351_),
    .Q(\cpu.regs[2][30] ));
 sg13g2_dfrbp_1 _12360_ (.CLK(net3799),
    .RESET_B(net107),
    .D(_00916_),
    .Q_N(_00350_),
    .Q(\cpu.regs[2][31] ));
 sg13g2_dfrbp_1 _12361_ (.CLK(net3752),
    .RESET_B(net106),
    .D(_00917_),
    .Q_N(_05998_),
    .Q(\irqvect[0][0] ));
 sg13g2_dfrbp_1 _12362_ (.CLK(net3753),
    .RESET_B(net105),
    .D(_00918_),
    .Q_N(_05997_),
    .Q(\irqvect[0][1] ));
 sg13g2_dfrbp_1 _12363_ (.CLK(net3751),
    .RESET_B(net104),
    .D(_00919_),
    .Q_N(_05996_),
    .Q(\irqvect[0][2] ));
 sg13g2_dfrbp_1 _12364_ (.CLK(net3755),
    .RESET_B(net103),
    .D(_00920_),
    .Q_N(_05995_),
    .Q(\irqvect[0][3] ));
 sg13g2_dfrbp_1 _12365_ (.CLK(net3755),
    .RESET_B(net102),
    .D(_00921_),
    .Q_N(_05994_),
    .Q(\irqvect[0][4] ));
 sg13g2_dfrbp_1 _12366_ (.CLK(net3753),
    .RESET_B(net101),
    .D(_00922_),
    .Q_N(_05993_),
    .Q(\irqvect[0][5] ));
 sg13g2_dfrbp_1 _12367_ (.CLK(net3754),
    .RESET_B(net100),
    .D(_00923_),
    .Q_N(_05992_),
    .Q(\irqvect[0][6] ));
 sg13g2_dfrbp_1 _12368_ (.CLK(net3754),
    .RESET_B(net99),
    .D(_00924_),
    .Q_N(_05991_),
    .Q(\irqvect[0][7] ));
 sg13g2_dfrbp_1 _12369_ (.CLK(net3760),
    .RESET_B(net98),
    .D(_00925_),
    .Q_N(_05990_),
    .Q(\irqvect[0][8] ));
 sg13g2_dfrbp_1 _12370_ (.CLK(net3746),
    .RESET_B(net97),
    .D(_00926_),
    .Q_N(_05989_),
    .Q(\irqvect[0][9] ));
 sg13g2_dfrbp_1 _12371_ (.CLK(net3756),
    .RESET_B(net96),
    .D(_00927_),
    .Q_N(_05988_),
    .Q(\irqvect[0][10] ));
 sg13g2_dfrbp_1 _12372_ (.CLK(net3742),
    .RESET_B(net95),
    .D(_00928_),
    .Q_N(_05987_),
    .Q(\irqvect[0][11] ));
 sg13g2_dfrbp_1 _12373_ (.CLK(net3745),
    .RESET_B(net94),
    .D(_00929_),
    .Q_N(_05986_),
    .Q(\irqvect[0][12] ));
 sg13g2_dfrbp_1 _12374_ (.CLK(net3758),
    .RESET_B(net93),
    .D(_00930_),
    .Q_N(_05985_),
    .Q(\irqvect[0][13] ));
 sg13g2_dfrbp_1 _12375_ (.CLK(net3750),
    .RESET_B(net92),
    .D(_00931_),
    .Q_N(_05984_),
    .Q(\irqvect[0][14] ));
 sg13g2_dfrbp_1 _12376_ (.CLK(net3751),
    .RESET_B(net91),
    .D(_00932_),
    .Q_N(_05983_),
    .Q(\irqvect[0][15] ));
 sg13g2_dfrbp_1 _12377_ (.CLK(net3750),
    .RESET_B(net90),
    .D(_00933_),
    .Q_N(_05982_),
    .Q(\irqvect[0][16] ));
 sg13g2_dfrbp_1 _12378_ (.CLK(net3745),
    .RESET_B(net89),
    .D(_00934_),
    .Q_N(_05981_),
    .Q(\irqvect[0][17] ));
 sg13g2_dfrbp_1 _12379_ (.CLK(net3744),
    .RESET_B(net88),
    .D(_00935_),
    .Q_N(_05980_),
    .Q(\irqvect[0][18] ));
 sg13g2_dfrbp_1 _12380_ (.CLK(net3740),
    .RESET_B(net87),
    .D(_00936_),
    .Q_N(_05979_),
    .Q(\irqvect[0][19] ));
 sg13g2_dfrbp_1 _12381_ (.CLK(net3740),
    .RESET_B(net86),
    .D(_00937_),
    .Q_N(_05978_),
    .Q(\irqvect[0][20] ));
 sg13g2_dfrbp_1 _12382_ (.CLK(net3746),
    .RESET_B(net85),
    .D(_00938_),
    .Q_N(_05977_),
    .Q(\irqvect[0][21] ));
 sg13g2_dfrbp_1 _12383_ (.CLK(net3743),
    .RESET_B(net84),
    .D(_00939_),
    .Q_N(_05976_),
    .Q(\irqvect[0][22] ));
 sg13g2_dfrbp_1 _12384_ (.CLK(net3743),
    .RESET_B(net83),
    .D(_00940_),
    .Q_N(_05975_),
    .Q(\irqvect[0][23] ));
 sg13g2_dfrbp_1 _12385_ (.CLK(net3743),
    .RESET_B(net82),
    .D(_00941_),
    .Q_N(_05974_),
    .Q(\irqvect[0][24] ));
 sg13g2_dfrbp_1 _12386_ (.CLK(net3756),
    .RESET_B(net81),
    .D(_00942_),
    .Q_N(_05973_),
    .Q(\irqvect[0][25] ));
 sg13g2_dfrbp_1 _12387_ (.CLK(net3744),
    .RESET_B(net80),
    .D(_00943_),
    .Q_N(_05972_),
    .Q(\irqvect[0][26] ));
 sg13g2_dfrbp_1 _12388_ (.CLK(net3747),
    .RESET_B(net79),
    .D(_00944_),
    .Q_N(_05971_),
    .Q(\irqvect[0][27] ));
 sg13g2_dfrbp_1 _12389_ (.CLK(net3741),
    .RESET_B(net78),
    .D(_00945_),
    .Q_N(_05970_),
    .Q(\irqvect[0][28] ));
 sg13g2_dfrbp_1 _12390_ (.CLK(net3741),
    .RESET_B(net77),
    .D(_00946_),
    .Q_N(_05969_),
    .Q(\irqvect[0][29] ));
 sg13g2_dfrbp_1 _12391_ (.CLK(net3840),
    .RESET_B(net76),
    .D(_00947_),
    .Q_N(_00349_),
    .Q(\cpu.regs[10][0] ));
 sg13g2_dfrbp_1 _12392_ (.CLK(net3844),
    .RESET_B(net75),
    .D(_00948_),
    .Q_N(_00348_),
    .Q(\cpu.regs[10][1] ));
 sg13g2_dfrbp_1 _12393_ (.CLK(net3795),
    .RESET_B(net74),
    .D(_00949_),
    .Q_N(_00347_),
    .Q(\cpu.regs[10][2] ));
 sg13g2_dfrbp_1 _12394_ (.CLK(net3862),
    .RESET_B(net73),
    .D(_00950_),
    .Q_N(_00346_),
    .Q(\cpu.regs[10][3] ));
 sg13g2_dfrbp_1 _12395_ (.CLK(net3844),
    .RESET_B(net72),
    .D(_00951_),
    .Q_N(_00345_),
    .Q(\cpu.regs[10][4] ));
 sg13g2_dfrbp_1 _12396_ (.CLK(net3864),
    .RESET_B(net71),
    .D(_00952_),
    .Q_N(_00344_),
    .Q(\cpu.regs[10][5] ));
 sg13g2_dfrbp_1 _12397_ (.CLK(net3847),
    .RESET_B(net70),
    .D(_00953_),
    .Q_N(_00343_),
    .Q(\cpu.regs[10][6] ));
 sg13g2_dfrbp_1 _12398_ (.CLK(net3864),
    .RESET_B(net69),
    .D(_00954_),
    .Q_N(_00342_),
    .Q(\cpu.regs[10][7] ));
 sg13g2_dfrbp_1 _12399_ (.CLK(net3868),
    .RESET_B(net68),
    .D(_00955_),
    .Q_N(_00341_),
    .Q(\cpu.regs[10][8] ));
 sg13g2_dfrbp_1 _12400_ (.CLK(net3845),
    .RESET_B(net67),
    .D(_00956_),
    .Q_N(_00340_),
    .Q(\cpu.regs[10][9] ));
 sg13g2_dfrbp_1 _12401_ (.CLK(net3858),
    .RESET_B(net66),
    .D(_00957_),
    .Q_N(_00339_),
    .Q(\cpu.regs[10][10] ));
 sg13g2_dfrbp_1 _12402_ (.CLK(net3857),
    .RESET_B(net65),
    .D(_00958_),
    .Q_N(_00338_),
    .Q(\cpu.regs[10][11] ));
 sg13g2_dfrbp_1 _12403_ (.CLK(net3807),
    .RESET_B(net64),
    .D(_00959_),
    .Q_N(_00337_),
    .Q(\cpu.regs[10][12] ));
 sg13g2_dfrbp_1 _12404_ (.CLK(net3806),
    .RESET_B(net63),
    .D(_00960_),
    .Q_N(_00336_),
    .Q(\cpu.regs[10][13] ));
 sg13g2_dfrbp_1 _12405_ (.CLK(net3854),
    .RESET_B(net62),
    .D(_00961_),
    .Q_N(_00335_),
    .Q(\cpu.regs[10][14] ));
 sg13g2_dfrbp_1 _12406_ (.CLK(net3851),
    .RESET_B(net61),
    .D(_00962_),
    .Q_N(_00334_),
    .Q(\cpu.regs[10][15] ));
 sg13g2_dfrbp_1 _12407_ (.CLK(net3837),
    .RESET_B(net60),
    .D(_00963_),
    .Q_N(_00333_),
    .Q(\cpu.regs[10][16] ));
 sg13g2_dfrbp_1 _12408_ (.CLK(net3859),
    .RESET_B(net59),
    .D(_00964_),
    .Q_N(_00332_),
    .Q(\cpu.regs[10][17] ));
 sg13g2_dfrbp_1 _12409_ (.CLK(net3832),
    .RESET_B(net58),
    .D(_00965_),
    .Q_N(_00331_),
    .Q(\cpu.regs[10][18] ));
 sg13g2_dfrbp_1 _12410_ (.CLK(net3830),
    .RESET_B(net57),
    .D(_00966_),
    .Q_N(_00330_),
    .Q(\cpu.regs[10][19] ));
 sg13g2_dfrbp_1 _12411_ (.CLK(net3803),
    .RESET_B(net56),
    .D(_00967_),
    .Q_N(_00329_),
    .Q(\cpu.regs[10][20] ));
 sg13g2_dfrbp_1 _12412_ (.CLK(net3819),
    .RESET_B(net55),
    .D(_00968_),
    .Q_N(_00328_),
    .Q(\cpu.regs[10][21] ));
 sg13g2_dfrbp_1 _12413_ (.CLK(net3814),
    .RESET_B(net54),
    .D(_00969_),
    .Q_N(_00327_),
    .Q(\cpu.regs[10][22] ));
 sg13g2_dfrbp_1 _12414_ (.CLK(net3818),
    .RESET_B(net53),
    .D(_00970_),
    .Q_N(_00326_),
    .Q(\cpu.regs[10][23] ));
 sg13g2_dfrbp_1 _12415_ (.CLK(net3813),
    .RESET_B(net52),
    .D(_00971_),
    .Q_N(_00325_),
    .Q(\cpu.regs[10][24] ));
 sg13g2_dfrbp_1 _12416_ (.CLK(net3822),
    .RESET_B(net51),
    .D(_00972_),
    .Q_N(_00324_),
    .Q(\cpu.regs[10][25] ));
 sg13g2_dfrbp_1 _12417_ (.CLK(net3804),
    .RESET_B(net50),
    .D(_00973_),
    .Q_N(_00323_),
    .Q(\cpu.regs[10][26] ));
 sg13g2_dfrbp_1 _12418_ (.CLK(net3817),
    .RESET_B(net49),
    .D(_00974_),
    .Q_N(_00322_),
    .Q(\cpu.regs[10][27] ));
 sg13g2_dfrbp_1 _12419_ (.CLK(net3824),
    .RESET_B(net48),
    .D(_00975_),
    .Q_N(_00321_),
    .Q(\cpu.regs[10][28] ));
 sg13g2_dfrbp_1 _12420_ (.CLK(net3826),
    .RESET_B(net47),
    .D(_00976_),
    .Q_N(_00320_),
    .Q(\cpu.regs[10][29] ));
 sg13g2_dfrbp_1 _12421_ (.CLK(net3809),
    .RESET_B(net46),
    .D(_00977_),
    .Q_N(_00319_),
    .Q(\cpu.regs[10][30] ));
 sg13g2_dfrbp_1 _12422_ (.CLK(net3802),
    .RESET_B(net45),
    .D(_00978_),
    .Q_N(_00318_),
    .Q(\cpu.regs[10][31] ));
 sg13g2_dfrbp_1 _12423_ (.CLK(net3750),
    .RESET_B(net44),
    .D(_00979_),
    .Q_N(_05968_),
    .Q(\irqvect[2][0] ));
 sg13g2_dfrbp_1 _12424_ (.CLK(net3753),
    .RESET_B(net43),
    .D(_00980_),
    .Q_N(_05967_),
    .Q(\irqvect[2][1] ));
 sg13g2_dfrbp_1 _12425_ (.CLK(net3751),
    .RESET_B(net42),
    .D(_00981_),
    .Q_N(_05966_),
    .Q(\irqvect[2][2] ));
 sg13g2_dfrbp_1 _12426_ (.CLK(net3755),
    .RESET_B(net41),
    .D(_00982_),
    .Q_N(_05965_),
    .Q(\irqvect[2][3] ));
 sg13g2_dfrbp_1 _12427_ (.CLK(net3779),
    .RESET_B(net40),
    .D(_00983_),
    .Q_N(_05964_),
    .Q(\irqvect[2][4] ));
 sg13g2_dfrbp_1 _12428_ (.CLK(net3754),
    .RESET_B(net39),
    .D(_00984_),
    .Q_N(_05963_),
    .Q(\irqvect[2][5] ));
 sg13g2_dfrbp_1 _12429_ (.CLK(net3754),
    .RESET_B(net38),
    .D(_00985_),
    .Q_N(_05962_),
    .Q(\irqvect[2][6] ));
 sg13g2_dfrbp_1 _12430_ (.CLK(net3755),
    .RESET_B(net37),
    .D(_00986_),
    .Q_N(_05961_),
    .Q(\irqvect[2][7] ));
 sg13g2_dfrbp_1 _12431_ (.CLK(net3759),
    .RESET_B(net36),
    .D(_00987_),
    .Q_N(_05960_),
    .Q(\irqvect[2][8] ));
 sg13g2_dfrbp_1 _12432_ (.CLK(net3746),
    .RESET_B(net35),
    .D(_00988_),
    .Q_N(_05959_),
    .Q(\irqvect[2][9] ));
 sg13g2_dfrbp_1 _12433_ (.CLK(net3751),
    .RESET_B(net34),
    .D(_00989_),
    .Q_N(_05958_),
    .Q(\irqvect[2][10] ));
 sg13g2_dfrbp_1 _12434_ (.CLK(net3742),
    .RESET_B(net33),
    .D(_00990_),
    .Q_N(_05957_),
    .Q(\irqvect[2][11] ));
 sg13g2_dfrbp_1 _12435_ (.CLK(net3747),
    .RESET_B(net32),
    .D(_00991_),
    .Q_N(_05956_),
    .Q(\irqvect[2][12] ));
 sg13g2_dfrbp_1 _12436_ (.CLK(net3758),
    .RESET_B(net31),
    .D(_00992_),
    .Q_N(_05955_),
    .Q(\irqvect[2][13] ));
 sg13g2_dfrbp_1 _12437_ (.CLK(net3752),
    .RESET_B(net30),
    .D(_00993_),
    .Q_N(_05954_),
    .Q(\irqvect[2][14] ));
 sg13g2_dfrbp_1 _12438_ (.CLK(net3751),
    .RESET_B(net29),
    .D(_00994_),
    .Q_N(_05953_),
    .Q(\irqvect[2][15] ));
 sg13g2_dfrbp_1 _12439_ (.CLK(net3750),
    .RESET_B(net28),
    .D(_00995_),
    .Q_N(_05952_),
    .Q(\irqvect[2][16] ));
 sg13g2_dfrbp_1 _12440_ (.CLK(net3745),
    .RESET_B(net27),
    .D(_00996_),
    .Q_N(_05951_),
    .Q(\irqvect[2][17] ));
 sg13g2_dfrbp_1 _12441_ (.CLK(net3744),
    .RESET_B(net26),
    .D(_00997_),
    .Q_N(_05950_),
    .Q(\irqvect[2][18] ));
 sg13g2_dfrbp_1 _12442_ (.CLK(net3740),
    .RESET_B(net25),
    .D(_00998_),
    .Q_N(_05949_),
    .Q(\irqvect[2][19] ));
 sg13g2_dfrbp_1 _12443_ (.CLK(net3740),
    .RESET_B(net24),
    .D(_00999_),
    .Q_N(_05948_),
    .Q(\irqvect[2][20] ));
 sg13g2_dfrbp_1 _12444_ (.CLK(net3746),
    .RESET_B(net23),
    .D(_01000_),
    .Q_N(_05947_),
    .Q(\irqvect[2][21] ));
 sg13g2_dfrbp_1 _12445_ (.CLK(net3748),
    .RESET_B(net22),
    .D(_01001_),
    .Q_N(_05946_),
    .Q(\irqvect[2][22] ));
 sg13g2_dfrbp_1 _12446_ (.CLK(net3743),
    .RESET_B(net21),
    .D(_01002_),
    .Q_N(_05945_),
    .Q(\irqvect[2][23] ));
 sg13g2_dfrbp_1 _12447_ (.CLK(net3743),
    .RESET_B(net20),
    .D(_01003_),
    .Q_N(_05944_),
    .Q(\irqvect[2][24] ));
 sg13g2_dfrbp_1 _12448_ (.CLK(net3757),
    .RESET_B(net19),
    .D(_01004_),
    .Q_N(_05943_),
    .Q(\irqvect[2][25] ));
 sg13g2_dfrbp_1 _12449_ (.CLK(net3744),
    .RESET_B(net18),
    .D(_01005_),
    .Q_N(_05942_),
    .Q(\irqvect[2][26] ));
 sg13g2_dfrbp_1 _12450_ (.CLK(net3756),
    .RESET_B(net17),
    .D(_01006_),
    .Q_N(_05941_),
    .Q(\irqvect[2][27] ));
 sg13g2_dfrbp_1 _12451_ (.CLK(net3740),
    .RESET_B(net889),
    .D(_01007_),
    .Q_N(_05940_),
    .Q(\irqvect[2][28] ));
 sg13g2_dfrbp_1 _12452_ (.CLK(net3741),
    .RESET_B(net888),
    .D(_01008_),
    .Q_N(_05939_),
    .Q(\irqvect[2][29] ));
 sg13g2_dfrbp_1 _12453_ (.CLK(net3840),
    .RESET_B(net887),
    .D(_01009_),
    .Q_N(_00317_),
    .Q(\cpu.regs[14][0] ));
 sg13g2_dfrbp_1 _12454_ (.CLK(net3841),
    .RESET_B(net886),
    .D(_01010_),
    .Q_N(_00316_),
    .Q(\cpu.regs[14][1] ));
 sg13g2_dfrbp_1 _12455_ (.CLK(net3793),
    .RESET_B(net885),
    .D(_01011_),
    .Q_N(_00315_),
    .Q(\cpu.regs[14][2] ));
 sg13g2_dfrbp_1 _12456_ (.CLK(net3855),
    .RESET_B(net884),
    .D(_01012_),
    .Q_N(_00314_),
    .Q(\cpu.regs[14][3] ));
 sg13g2_dfrbp_1 _12457_ (.CLK(net3793),
    .RESET_B(net883),
    .D(_01013_),
    .Q_N(_00313_),
    .Q(\cpu.regs[14][4] ));
 sg13g2_dfrbp_1 _12458_ (.CLK(net3867),
    .RESET_B(net882),
    .D(_01014_),
    .Q_N(_00312_),
    .Q(\cpu.regs[14][5] ));
 sg13g2_dfrbp_1 _12459_ (.CLK(net3846),
    .RESET_B(net881),
    .D(_01015_),
    .Q_N(_00311_),
    .Q(\cpu.regs[14][6] ));
 sg13g2_dfrbp_1 _12460_ (.CLK(net3861),
    .RESET_B(net880),
    .D(_01016_),
    .Q_N(_00310_),
    .Q(\cpu.regs[14][7] ));
 sg13g2_dfrbp_1 _12461_ (.CLK(net3866),
    .RESET_B(net879),
    .D(_01017_),
    .Q_N(_00309_),
    .Q(\cpu.regs[14][8] ));
 sg13g2_dfrbp_1 _12462_ (.CLK(net3862),
    .RESET_B(net878),
    .D(_01018_),
    .Q_N(_00308_),
    .Q(\cpu.regs[14][9] ));
 sg13g2_dfrbp_1 _12463_ (.CLK(net3868),
    .RESET_B(net877),
    .D(_01019_),
    .Q_N(_00307_),
    .Q(\cpu.regs[14][10] ));
 sg13g2_dfrbp_1 _12464_ (.CLK(net3857),
    .RESET_B(net876),
    .D(_01020_),
    .Q_N(_00306_),
    .Q(\cpu.regs[14][11] ));
 sg13g2_dfrbp_1 _12465_ (.CLK(net3804),
    .RESET_B(net875),
    .D(_01021_),
    .Q_N(_00305_),
    .Q(\cpu.regs[14][12] ));
 sg13g2_dfrbp_1 _12466_ (.CLK(net3806),
    .RESET_B(net874),
    .D(_01022_),
    .Q_N(_00304_),
    .Q(\cpu.regs[14][13] ));
 sg13g2_dfrbp_1 _12467_ (.CLK(net3854),
    .RESET_B(net873),
    .D(_01023_),
    .Q_N(_00303_),
    .Q(\cpu.regs[14][14] ));
 sg13g2_dfrbp_1 _12468_ (.CLK(net3852),
    .RESET_B(net872),
    .D(_01024_),
    .Q_N(_00302_),
    .Q(\cpu.regs[14][15] ));
 sg13g2_dfrbp_1 _12469_ (.CLK(net3837),
    .RESET_B(net871),
    .D(_01025_),
    .Q_N(_00301_),
    .Q(\cpu.regs[14][16] ));
 sg13g2_dfrbp_1 _12470_ (.CLK(net3858),
    .RESET_B(net870),
    .D(_01026_),
    .Q_N(_00300_),
    .Q(\cpu.regs[14][17] ));
 sg13g2_dfrbp_1 _12471_ (.CLK(net3829),
    .RESET_B(net869),
    .D(_01027_),
    .Q_N(_00299_),
    .Q(\cpu.regs[14][18] ));
 sg13g2_dfrbp_1 _12472_ (.CLK(net3830),
    .RESET_B(net868),
    .D(_01028_),
    .Q_N(_00298_),
    .Q(\cpu.regs[14][19] ));
 sg13g2_dfrbp_1 _12473_ (.CLK(net3803),
    .RESET_B(net867),
    .D(_01029_),
    .Q_N(_00297_),
    .Q(\cpu.regs[14][20] ));
 sg13g2_dfrbp_1 _12474_ (.CLK(net3821),
    .RESET_B(net866),
    .D(_01030_),
    .Q_N(_00296_),
    .Q(\cpu.regs[14][21] ));
 sg13g2_dfrbp_1 _12475_ (.CLK(net3815),
    .RESET_B(net865),
    .D(_01031_),
    .Q_N(_00295_),
    .Q(\cpu.regs[14][22] ));
 sg13g2_dfrbp_1 _12476_ (.CLK(net3816),
    .RESET_B(net864),
    .D(_01032_),
    .Q_N(_00294_),
    .Q(\cpu.regs[14][23] ));
 sg13g2_dfrbp_1 _12477_ (.CLK(net3816),
    .RESET_B(net863),
    .D(_01033_),
    .Q_N(_00293_),
    .Q(\cpu.regs[14][24] ));
 sg13g2_dfrbp_1 _12478_ (.CLK(net3829),
    .RESET_B(net862),
    .D(_01034_),
    .Q_N(_00292_),
    .Q(\cpu.regs[14][25] ));
 sg13g2_dfrbp_1 _12479_ (.CLK(net3813),
    .RESET_B(net861),
    .D(_01035_),
    .Q_N(_00291_),
    .Q(\cpu.regs[14][26] ));
 sg13g2_dfrbp_1 _12480_ (.CLK(net3825),
    .RESET_B(net860),
    .D(_01036_),
    .Q_N(_00290_),
    .Q(\cpu.regs[14][27] ));
 sg13g2_dfrbp_1 _12481_ (.CLK(net3817),
    .RESET_B(net859),
    .D(_01037_),
    .Q_N(_00289_),
    .Q(\cpu.regs[14][28] ));
 sg13g2_dfrbp_1 _12482_ (.CLK(net3826),
    .RESET_B(net858),
    .D(_01038_),
    .Q_N(_00288_),
    .Q(\cpu.regs[14][29] ));
 sg13g2_dfrbp_1 _12483_ (.CLK(net3809),
    .RESET_B(net857),
    .D(_01039_),
    .Q_N(_00287_),
    .Q(\cpu.regs[14][30] ));
 sg13g2_dfrbp_1 _12484_ (.CLK(net3813),
    .RESET_B(net856),
    .D(_01040_),
    .Q_N(_00286_),
    .Q(\cpu.regs[14][31] ));
 sg13g2_dfrbp_1 _12485_ (.CLK(net3794),
    .RESET_B(net855),
    .D(_01041_),
    .Q_N(_00285_),
    .Q(\cpu.regs[6][0] ));
 sg13g2_dfrbp_1 _12486_ (.CLK(net3842),
    .RESET_B(net854),
    .D(_01042_),
    .Q_N(_00284_),
    .Q(\cpu.regs[6][1] ));
 sg13g2_dfrbp_1 _12487_ (.CLK(net3793),
    .RESET_B(net853),
    .D(_01043_),
    .Q_N(_00283_),
    .Q(\cpu.regs[6][2] ));
 sg13g2_dfrbp_1 _12488_ (.CLK(net3846),
    .RESET_B(net852),
    .D(_01044_),
    .Q_N(_00282_),
    .Q(\cpu.regs[6][3] ));
 sg13g2_dfrbp_1 _12489_ (.CLK(net3789),
    .RESET_B(net851),
    .D(_01045_),
    .Q_N(_00281_),
    .Q(\cpu.regs[6][4] ));
 sg13g2_dfrbp_1 _12490_ (.CLK(net3863),
    .RESET_B(net850),
    .D(_01046_),
    .Q_N(_00280_),
    .Q(\cpu.regs[6][5] ));
 sg13g2_dfrbp_1 _12491_ (.CLK(net3843),
    .RESET_B(net849),
    .D(_01047_),
    .Q_N(_00279_),
    .Q(\cpu.regs[6][6] ));
 sg13g2_dfrbp_1 _12492_ (.CLK(net3848),
    .RESET_B(net848),
    .D(_01048_),
    .Q_N(_00278_),
    .Q(\cpu.regs[6][7] ));
 sg13g2_dfrbp_1 _12493_ (.CLK(net3862),
    .RESET_B(net847),
    .D(_01049_),
    .Q_N(_00277_),
    .Q(\cpu.regs[6][8] ));
 sg13g2_dfrbp_1 _12494_ (.CLK(net3834),
    .RESET_B(net846),
    .D(_01050_),
    .Q_N(_00276_),
    .Q(\cpu.regs[6][9] ));
 sg13g2_dfrbp_1 _12495_ (.CLK(net3853),
    .RESET_B(net845),
    .D(_01051_),
    .Q_N(_00275_),
    .Q(\cpu.regs[6][10] ));
 sg13g2_dfrbp_1 _12496_ (.CLK(net3856),
    .RESET_B(net844),
    .D(_01052_),
    .Q_N(_00274_),
    .Q(\cpu.regs[6][11] ));
 sg13g2_dfrbp_1 _12497_ (.CLK(net3761),
    .RESET_B(net843),
    .D(_01053_),
    .Q_N(_00273_),
    .Q(\cpu.regs[6][12] ));
 sg13g2_dfrbp_1 _12498_ (.CLK(net3761),
    .RESET_B(net842),
    .D(_01054_),
    .Q_N(_00272_),
    .Q(\cpu.regs[6][13] ));
 sg13g2_dfrbp_1 _12499_ (.CLK(net3836),
    .RESET_B(net841),
    .D(_01055_),
    .Q_N(_00271_),
    .Q(\cpu.regs[6][14] ));
 sg13g2_dfrbp_1 _12500_ (.CLK(net3835),
    .RESET_B(net840),
    .D(_01056_),
    .Q_N(_00270_),
    .Q(\cpu.regs[6][15] ));
 sg13g2_dfrbp_1 _12501_ (.CLK(net3841),
    .RESET_B(net839),
    .D(_01057_),
    .Q_N(_00269_),
    .Q(\cpu.regs[6][16] ));
 sg13g2_dfrbp_1 _12502_ (.CLK(net3853),
    .RESET_B(net838),
    .D(_01058_),
    .Q_N(_00268_),
    .Q(\cpu.regs[6][17] ));
 sg13g2_dfrbp_1 _12503_ (.CLK(net3831),
    .RESET_B(net837),
    .D(_01059_),
    .Q_N(_00267_),
    .Q(\cpu.regs[6][18] ));
 sg13g2_dfrbp_1 _12504_ (.CLK(net3852),
    .RESET_B(net836),
    .D(_01060_),
    .Q_N(_00266_),
    .Q(\cpu.regs[6][19] ));
 sg13g2_dfrbp_1 _12505_ (.CLK(net3761),
    .RESET_B(net835),
    .D(_01061_),
    .Q_N(_00265_),
    .Q(\cpu.regs[6][20] ));
 sg13g2_dfrbp_1 _12506_ (.CLK(net3822),
    .RESET_B(net834),
    .D(_01062_),
    .Q_N(_00264_),
    .Q(\cpu.regs[6][21] ));
 sg13g2_dfrbp_1 _12507_ (.CLK(net3829),
    .RESET_B(net833),
    .D(_01063_),
    .Q_N(_00263_),
    .Q(\cpu.regs[6][22] ));
 sg13g2_dfrbp_1 _12508_ (.CLK(net3820),
    .RESET_B(net832),
    .D(_01064_),
    .Q_N(_00262_),
    .Q(\cpu.regs[6][23] ));
 sg13g2_dfrbp_1 _12509_ (.CLK(net3806),
    .RESET_B(net831),
    .D(_01065_),
    .Q_N(_00261_),
    .Q(\cpu.regs[6][24] ));
 sg13g2_dfrbp_1 _12510_ (.CLK(net3822),
    .RESET_B(net830),
    .D(_01066_),
    .Q_N(_00260_),
    .Q(\cpu.regs[6][25] ));
 sg13g2_dfrbp_1 _12511_ (.CLK(net3800),
    .RESET_B(net829),
    .D(_01067_),
    .Q_N(_00259_),
    .Q(\cpu.regs[6][26] ));
 sg13g2_dfrbp_1 _12512_ (.CLK(net3824),
    .RESET_B(net828),
    .D(_01068_),
    .Q_N(_00258_),
    .Q(\cpu.regs[6][27] ));
 sg13g2_dfrbp_1 _12513_ (.CLK(net3809),
    .RESET_B(net827),
    .D(_01069_),
    .Q_N(_00257_),
    .Q(\cpu.regs[6][28] ));
 sg13g2_dfrbp_1 _12514_ (.CLK(net3827),
    .RESET_B(net826),
    .D(_01070_),
    .Q_N(_00256_),
    .Q(\cpu.regs[6][29] ));
 sg13g2_dfrbp_1 _12515_ (.CLK(net3763),
    .RESET_B(net825),
    .D(_01071_),
    .Q_N(_00255_),
    .Q(\cpu.regs[6][30] ));
 sg13g2_dfrbp_1 _12516_ (.CLK(net3768),
    .RESET_B(net824),
    .D(_01072_),
    .Q_N(_00254_),
    .Q(\cpu.regs[6][31] ));
 sg13g2_dfrbp_1 _12517_ (.CLK(net3794),
    .RESET_B(net823),
    .D(_01073_),
    .Q_N(_00253_),
    .Q(\cpu.regs[5][0] ));
 sg13g2_dfrbp_1 _12518_ (.CLK(net3842),
    .RESET_B(net822),
    .D(_01074_),
    .Q_N(_00252_),
    .Q(\cpu.regs[5][1] ));
 sg13g2_dfrbp_1 _12519_ (.CLK(net3792),
    .RESET_B(net821),
    .D(_01075_),
    .Q_N(_00251_),
    .Q(\cpu.regs[5][2] ));
 sg13g2_dfrbp_1 _12520_ (.CLK(net3846),
    .RESET_B(net820),
    .D(_01076_),
    .Q_N(_00250_),
    .Q(\cpu.regs[5][3] ));
 sg13g2_dfrbp_1 _12521_ (.CLK(net3789),
    .RESET_B(net819),
    .D(_01077_),
    .Q_N(_00249_),
    .Q(\cpu.regs[5][4] ));
 sg13g2_dfrbp_1 _12522_ (.CLK(net3865),
    .RESET_B(net787),
    .D(_01078_),
    .Q_N(_00248_),
    .Q(\cpu.regs[5][5] ));
 sg13g2_dfrbp_1 _12523_ (.CLK(net3843),
    .RESET_B(net786),
    .D(_01079_),
    .Q_N(_00247_),
    .Q(\cpu.regs[5][6] ));
 sg13g2_dfrbp_1 _12524_ (.CLK(net3848),
    .RESET_B(net785),
    .D(_01080_),
    .Q_N(_00246_),
    .Q(\cpu.regs[5][7] ));
 sg13g2_dfrbp_1 _12525_ (.CLK(net3845),
    .RESET_B(net784),
    .D(_01081_),
    .Q_N(_00245_),
    .Q(\cpu.regs[5][8] ));
 sg13g2_dfrbp_1 _12526_ (.CLK(net3834),
    .RESET_B(net783),
    .D(_01082_),
    .Q_N(_00244_),
    .Q(\cpu.regs[5][9] ));
 sg13g2_dfrbp_1 _12527_ (.CLK(net3861),
    .RESET_B(net782),
    .D(_01083_),
    .Q_N(_00243_),
    .Q(\cpu.regs[5][10] ));
 sg13g2_dfrbp_1 _12528_ (.CLK(net3852),
    .RESET_B(net781),
    .D(_01084_),
    .Q_N(_00242_),
    .Q(\cpu.regs[5][11] ));
 sg13g2_dfrbp_1 _12529_ (.CLK(net3761),
    .RESET_B(net780),
    .D(_01085_),
    .Q_N(_00241_),
    .Q(\cpu.regs[5][12] ));
 sg13g2_dfrbp_1 _12530_ (.CLK(net3762),
    .RESET_B(net779),
    .D(_01086_),
    .Q_N(_00240_),
    .Q(\cpu.regs[5][13] ));
 sg13g2_dfrbp_1 _12531_ (.CLK(net3834),
    .RESET_B(net778),
    .D(_01087_),
    .Q_N(_00239_),
    .Q(\cpu.regs[5][14] ));
 sg13g2_dfrbp_1 _12532_ (.CLK(net3835),
    .RESET_B(net777),
    .D(_01088_),
    .Q_N(_00238_),
    .Q(\cpu.regs[5][15] ));
 sg13g2_dfrbp_1 _12533_ (.CLK(net3839),
    .RESET_B(net776),
    .D(_01089_),
    .Q_N(_00237_),
    .Q(\cpu.regs[5][16] ));
 sg13g2_dfrbp_1 _12534_ (.CLK(net3853),
    .RESET_B(net775),
    .D(_01090_),
    .Q_N(_00236_),
    .Q(\cpu.regs[5][17] ));
 sg13g2_dfrbp_1 _12535_ (.CLK(net3831),
    .RESET_B(net774),
    .D(_01091_),
    .Q_N(_00235_),
    .Q(\cpu.regs[5][18] ));
 sg13g2_dfrbp_1 _12536_ (.CLK(net3826),
    .RESET_B(net773),
    .D(_01092_),
    .Q_N(_00234_),
    .Q(\cpu.regs[5][19] ));
 sg13g2_dfrbp_1 _12537_ (.CLK(net3762),
    .RESET_B(net772),
    .D(_01093_),
    .Q_N(_00233_),
    .Q(\cpu.regs[5][20] ));
 sg13g2_dfrbp_1 _12538_ (.CLK(net3818),
    .RESET_B(net771),
    .D(_01094_),
    .Q_N(_00232_),
    .Q(\cpu.regs[5][21] ));
 sg13g2_dfrbp_1 _12539_ (.CLK(net3824),
    .RESET_B(net770),
    .D(_01095_),
    .Q_N(_00231_),
    .Q(\cpu.regs[5][22] ));
 sg13g2_dfrbp_1 _12540_ (.CLK(net3820),
    .RESET_B(net769),
    .D(_01096_),
    .Q_N(_00230_),
    .Q(\cpu.regs[5][23] ));
 sg13g2_dfrbp_1 _12541_ (.CLK(net3806),
    .RESET_B(net768),
    .D(_01097_),
    .Q_N(_00229_),
    .Q(\cpu.regs[5][24] ));
 sg13g2_dfrbp_1 _12542_ (.CLK(net3821),
    .RESET_B(net767),
    .D(_01098_),
    .Q_N(_00228_),
    .Q(\cpu.regs[5][25] ));
 sg13g2_dfrbp_1 _12543_ (.CLK(net3801),
    .RESET_B(net766),
    .D(_01099_),
    .Q_N(_00227_),
    .Q(\cpu.regs[5][26] ));
 sg13g2_dfrbp_1 _12544_ (.CLK(net3824),
    .RESET_B(net765),
    .D(_01100_),
    .Q_N(_00226_),
    .Q(\cpu.regs[5][27] ));
 sg13g2_dfrbp_1 _12545_ (.CLK(net3810),
    .RESET_B(net764),
    .D(_01101_),
    .Q_N(_00225_),
    .Q(\cpu.regs[5][28] ));
 sg13g2_dfrbp_1 _12546_ (.CLK(net3811),
    .RESET_B(net763),
    .D(_01102_),
    .Q_N(_00224_),
    .Q(\cpu.regs[5][29] ));
 sg13g2_dfrbp_1 _12547_ (.CLK(net3763),
    .RESET_B(net762),
    .D(_01103_),
    .Q_N(_00223_),
    .Q(\cpu.regs[5][30] ));
 sg13g2_dfrbp_1 _12548_ (.CLK(net3767),
    .RESET_B(net761),
    .D(_01104_),
    .Q_N(_00222_),
    .Q(\cpu.regs[5][31] ));
 sg13g2_dfrbp_1 _12549_ (.CLK(net3919),
    .RESET_B(net3718),
    .D(_01105_),
    .Q_N(txd),
    .Q(_00572_));
 sg13g2_dfrbp_1 _12550_ (.CLK(net3919),
    .RESET_B(net3715),
    .D(_01106_),
    .Q_N(\uart0.txsh[1] ),
    .Q(_00573_));
 sg13g2_dfrbp_1 _12551_ (.CLK(net3919),
    .RESET_B(net3715),
    .D(_01107_),
    .Q_N(\uart0.txsh[2] ),
    .Q(_00574_));
 sg13g2_dfrbp_1 _12552_ (.CLK(net3917),
    .RESET_B(net3717),
    .D(_01108_),
    .Q_N(\uart0.txsh[3] ),
    .Q(_00575_));
 sg13g2_dfrbp_1 _12553_ (.CLK(net3917),
    .RESET_B(net3715),
    .D(_01109_),
    .Q_N(\uart0.txsh[4] ),
    .Q(_00576_));
 sg13g2_dfrbp_1 _12554_ (.CLK(net3919),
    .RESET_B(net3715),
    .D(_01110_),
    .Q_N(\uart0.txsh[5] ),
    .Q(_00577_));
 sg13g2_dfrbp_1 _12555_ (.CLK(net3917),
    .RESET_B(net3715),
    .D(_01111_),
    .Q_N(\uart0.txsh[6] ),
    .Q(_00578_));
 sg13g2_dfrbp_1 _12556_ (.CLK(net3917),
    .RESET_B(net3716),
    .D(_01112_),
    .Q_N(\uart0.txsh[7] ),
    .Q(_00579_));
 sg13g2_dfrbp_1 _12557_ (.CLK(net3917),
    .RESET_B(net3716),
    .D(_01113_),
    .Q_N(\uart0.txsh[8] ),
    .Q(_00580_));
 sg13g2_dfrbp_1 _12558_ (.CLK(net3790),
    .RESET_B(net3722),
    .D(_00004_),
    .Q_N(_06029_),
    .Q(\pwmc[0] ));
 sg13g2_dfrbp_1 _12559_ (.CLK(net3790),
    .RESET_B(net3721),
    .D(_00005_),
    .Q_N(_06030_),
    .Q(\pwmc[1] ));
 sg13g2_dfrbp_1 _12560_ (.CLK(net3791),
    .RESET_B(net3720),
    .D(_00006_),
    .Q_N(_00542_),
    .Q(\pwmc[2] ));
 sg13g2_dfrbp_1 _12561_ (.CLK(net3790),
    .RESET_B(net3720),
    .D(_00007_),
    .Q_N(_06031_),
    .Q(\pwmc[3] ));
 sg13g2_dfrbp_1 _12562_ (.CLK(net3791),
    .RESET_B(net3720),
    .D(_00008_),
    .Q_N(_00543_),
    .Q(\pwmc[4] ));
 sg13g2_dfrbp_1 _12563_ (.CLK(net3789),
    .RESET_B(net3720),
    .D(_00009_),
    .Q_N(_06032_),
    .Q(\pwmc[5] ));
 sg13g2_dfrbp_1 _12564_ (.CLK(net3789),
    .RESET_B(net3720),
    .D(_00010_),
    .Q_N(_06033_),
    .Q(\pwmc[6] ));
 sg13g2_dfrbp_1 _12565_ (.CLK(net3791),
    .RESET_B(net3720),
    .D(_00011_),
    .Q_N(_05938_),
    .Q(\pwmc[7] ));
 sg13g2_dfrbp_1 _12566_ (.CLK(net3779),
    .RESET_B(net3719),
    .D(_01114_),
    .Q_N(_05937_),
    .Q(\irqen[0] ));
 sg13g2_dfrbp_1 _12567_ (.CLK(net3779),
    .RESET_B(net3719),
    .D(_01115_),
    .Q_N(_05936_),
    .Q(\irqen[1] ));
 sg13g2_dfrbp_1 _12568_ (.CLK(net3780),
    .RESET_B(net3717),
    .D(_01116_),
    .Q_N(_05935_),
    .Q(\irqen[2] ));
 sg13g2_dfrbp_1 _12569_ (.CLK(net3779),
    .RESET_B(net3705),
    .D(_01117_),
    .Q_N(_05934_),
    .Q(\irqen[3] ));
 sg13g2_dfrbp_1 _12570_ (.CLK(net3779),
    .RESET_B(net3717),
    .D(_01118_),
    .Q_N(_05933_),
    .Q(\irqen[4] ));
 sg13g2_dfrbp_1 _12571_ (.CLK(net3789),
    .RESET_B(net701),
    .D(_01119_),
    .Q_N(_05932_),
    .Q(\pwmbuf[0] ));
 sg13g2_dfrbp_1 _12572_ (.CLK(net3787),
    .RESET_B(net700),
    .D(_01120_),
    .Q_N(_05931_),
    .Q(\pwmbuf[1] ));
 sg13g2_dfrbp_1 _12573_ (.CLK(net3787),
    .RESET_B(net699),
    .D(_01121_),
    .Q_N(_05930_),
    .Q(\pwmbuf[2] ));
 sg13g2_dfrbp_1 _12574_ (.CLK(net3789),
    .RESET_B(net698),
    .D(_01122_),
    .Q_N(_05929_),
    .Q(\pwmbuf[3] ));
 sg13g2_dfrbp_1 _12575_ (.CLK(net3788),
    .RESET_B(net697),
    .D(_01123_),
    .Q_N(_05928_),
    .Q(\pwmbuf[4] ));
 sg13g2_dfrbp_1 _12576_ (.CLK(net3789),
    .RESET_B(net696),
    .D(_01124_),
    .Q_N(_05927_),
    .Q(\pwmbuf[5] ));
 sg13g2_dfrbp_1 _12577_ (.CLK(net3790),
    .RESET_B(net695),
    .D(_01125_),
    .Q_N(_05926_),
    .Q(\pwmbuf[6] ));
 sg13g2_dfrbp_1 _12578_ (.CLK(net3791),
    .RESET_B(net694),
    .D(_01126_),
    .Q_N(_05925_),
    .Q(\pwmbuf[7] ));
 sg13g2_dfrbp_1 _12579_ (.CLK(net3788),
    .RESET_B(net693),
    .D(_01127_),
    .Q_N(_05924_),
    .Q(\pwm[0] ));
 sg13g2_dfrbp_1 _12580_ (.CLK(net3787),
    .RESET_B(net692),
    .D(_01128_),
    .Q_N(_05923_),
    .Q(\pwm[1] ));
 sg13g2_dfrbp_1 _12581_ (.CLK(net3787),
    .RESET_B(net691),
    .D(_01129_),
    .Q_N(_05922_),
    .Q(\pwm[2] ));
 sg13g2_dfrbp_1 _12582_ (.CLK(net3787),
    .RESET_B(net690),
    .D(_01130_),
    .Q_N(_05921_),
    .Q(\pwm[3] ));
 sg13g2_dfrbp_1 _12583_ (.CLK(net3788),
    .RESET_B(net689),
    .D(_01131_),
    .Q_N(_05920_),
    .Q(\pwm[4] ));
 sg13g2_dfrbp_1 _12584_ (.CLK(net3787),
    .RESET_B(net688),
    .D(_01132_),
    .Q_N(_05919_),
    .Q(\pwm[5] ));
 sg13g2_dfrbp_1 _12585_ (.CLK(net3789),
    .RESET_B(net687),
    .D(_01133_),
    .Q_N(_05918_),
    .Q(\pwm[6] ));
 sg13g2_dfrbp_1 _12586_ (.CLK(net3791),
    .RESET_B(net686),
    .D(_01134_),
    .Q_N(_05917_),
    .Q(\pwm[7] ));
 sg13g2_dfrbp_1 _12587_ (.CLK(net3791),
    .RESET_B(net3720),
    .D(_01135_),
    .Q_N(_05916_),
    .Q(pwmout));
 sg13g2_dfrbp_1 _12588_ (.CLK(net3780),
    .RESET_B(net685),
    .D(_01136_),
    .Q_N(_05915_),
    .Q(udirty));
 sg13g2_dfrbp_1 _12589_ (.CLK(net3915),
    .RESET_B(net683),
    .D(_05639_),
    .Q_N(_05639_),
    .Q(\tcount[0] ));
 sg13g2_dfrbp_1 _12590_ (.CLK(net3918),
    .RESET_B(net682),
    .D(_00038_),
    .Q_N(_05914_),
    .Q(\tcount[1] ));
 sg13g2_dfrbp_1 _12591_ (.CLK(net3918),
    .RESET_B(net681),
    .D(_00049_),
    .Q_N(_05913_),
    .Q(\tcount[2] ));
 sg13g2_dfrbp_1 _12592_ (.CLK(net3914),
    .RESET_B(net680),
    .D(_00052_),
    .Q_N(_05912_),
    .Q(\tcount[3] ));
 sg13g2_dfrbp_1 _12593_ (.CLK(net3914),
    .RESET_B(net679),
    .D(_00053_),
    .Q_N(_05911_),
    .Q(\tcount[4] ));
 sg13g2_dfrbp_1 _12594_ (.CLK(net3918),
    .RESET_B(net678),
    .D(_00054_),
    .Q_N(_05910_),
    .Q(\tcount[5] ));
 sg13g2_dfrbp_1 _12595_ (.CLK(net3918),
    .RESET_B(net677),
    .D(_00055_),
    .Q_N(_05909_),
    .Q(\tcount[6] ));
 sg13g2_dfrbp_1 _12596_ (.CLK(net3918),
    .RESET_B(net676),
    .D(_00056_),
    .Q_N(_05908_),
    .Q(\tcount[7] ));
 sg13g2_dfrbp_1 _12597_ (.CLK(net3918),
    .RESET_B(net675),
    .D(_00057_),
    .Q_N(_05907_),
    .Q(\tcount[8] ));
 sg13g2_dfrbp_1 _12598_ (.CLK(net3918),
    .RESET_B(net674),
    .D(_00058_),
    .Q_N(_05906_),
    .Q(\tcount[9] ));
 sg13g2_dfrbp_1 _12599_ (.CLK(net3919),
    .RESET_B(net673),
    .D(_00028_),
    .Q_N(_05905_),
    .Q(\tcount[10] ));
 sg13g2_dfrbp_1 _12600_ (.CLK(net3923),
    .RESET_B(net672),
    .D(_00029_),
    .Q_N(_05904_),
    .Q(\tcount[11] ));
 sg13g2_dfrbp_1 _12601_ (.CLK(net3923),
    .RESET_B(net671),
    .D(_00030_),
    .Q_N(_05903_),
    .Q(\tcount[12] ));
 sg13g2_dfrbp_1 _12602_ (.CLK(net3921),
    .RESET_B(net670),
    .D(_00031_),
    .Q_N(_05902_),
    .Q(\tcount[13] ));
 sg13g2_dfrbp_1 _12603_ (.CLK(net3922),
    .RESET_B(net669),
    .D(_00032_),
    .Q_N(_05901_),
    .Q(\tcount[14] ));
 sg13g2_dfrbp_1 _12604_ (.CLK(net3921),
    .RESET_B(net668),
    .D(_00033_),
    .Q_N(_05900_),
    .Q(\tcount[15] ));
 sg13g2_dfrbp_1 _12605_ (.CLK(net3921),
    .RESET_B(net667),
    .D(_00034_),
    .Q_N(_05899_),
    .Q(\tcount[16] ));
 sg13g2_dfrbp_1 _12606_ (.CLK(net3921),
    .RESET_B(net666),
    .D(_00035_),
    .Q_N(_05898_),
    .Q(\tcount[17] ));
 sg13g2_dfrbp_1 _12607_ (.CLK(net3921),
    .RESET_B(net665),
    .D(_00036_),
    .Q_N(_05897_),
    .Q(\tcount[18] ));
 sg13g2_dfrbp_1 _12608_ (.CLK(net3921),
    .RESET_B(net664),
    .D(_00037_),
    .Q_N(_05896_),
    .Q(\tcount[19] ));
 sg13g2_dfrbp_1 _12609_ (.CLK(net3922),
    .RESET_B(net663),
    .D(_00039_),
    .Q_N(_05895_),
    .Q(\tcount[20] ));
 sg13g2_dfrbp_1 _12610_ (.CLK(net3922),
    .RESET_B(net662),
    .D(_00040_),
    .Q_N(_05894_),
    .Q(\tcount[21] ));
 sg13g2_dfrbp_1 _12611_ (.CLK(net3922),
    .RESET_B(net661),
    .D(_00041_),
    .Q_N(_05893_),
    .Q(\tcount[22] ));
 sg13g2_dfrbp_1 _12612_ (.CLK(net3922),
    .RESET_B(net660),
    .D(_00042_),
    .Q_N(_05892_),
    .Q(\tcount[23] ));
 sg13g2_dfrbp_1 _12613_ (.CLK(net3922),
    .RESET_B(net659),
    .D(_00043_),
    .Q_N(_05891_),
    .Q(\tcount[24] ));
 sg13g2_dfrbp_1 _12614_ (.CLK(net3924),
    .RESET_B(net658),
    .D(_00044_),
    .Q_N(_05890_),
    .Q(\tcount[25] ));
 sg13g2_dfrbp_1 _12615_ (.CLK(net3924),
    .RESET_B(net657),
    .D(_00045_),
    .Q_N(_05889_),
    .Q(\tcount[26] ));
 sg13g2_dfrbp_1 _12616_ (.CLK(net3923),
    .RESET_B(net656),
    .D(_00046_),
    .Q_N(_05888_),
    .Q(\tcount[27] ));
 sg13g2_dfrbp_1 _12617_ (.CLK(net3924),
    .RESET_B(net655),
    .D(_00047_),
    .Q_N(_05887_),
    .Q(\tcount[28] ));
 sg13g2_dfrbp_1 _12618_ (.CLK(net3923),
    .RESET_B(net654),
    .D(_00048_),
    .Q_N(_05886_),
    .Q(\tcount[29] ));
 sg13g2_dfrbp_1 _12619_ (.CLK(net3923),
    .RESET_B(net653),
    .D(_00050_),
    .Q_N(_05885_),
    .Q(\tcount[30] ));
 sg13g2_dfrbp_1 _12620_ (.CLK(net3923),
    .RESET_B(net652),
    .D(_00051_),
    .Q_N(_05884_),
    .Q(\tcount[31] ));
 sg13g2_dfrbp_1 _12621_ (.CLK(net3798),
    .RESET_B(net3719),
    .D(_01137_),
    .Q_N(_05883_),
    .Q(pwmirq));
 sg13g2_dfrbp_1 _12622_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net651),
    .D(_01138_),
    .Q_N(_05882_),
    .Q(\xdi[0] ));
 sg13g2_dfrbp_1 _12623_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net650),
    .D(net915),
    .Q_N(_05881_),
    .Q(\xdi[1] ));
 sg13g2_dfrbp_1 _12624_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net649),
    .D(net902),
    .Q_N(_05880_),
    .Q(\xdi[2] ));
 sg13g2_dfrbp_1 _12625_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net648),
    .D(_01141_),
    .Q_N(_05879_),
    .Q(\xdi[3] ));
 sg13g2_dfrbp_1 _12626_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net647),
    .D(_01142_),
    .Q_N(_05878_),
    .Q(\xdi[4] ));
 sg13g2_dfrbp_1 _12627_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net646),
    .D(net898),
    .Q_N(_05877_),
    .Q(\xdi[5] ));
 sg13g2_dfrbp_1 _12628_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net645),
    .D(_01144_),
    .Q_N(_05876_),
    .Q(\xdi[6] ));
 sg13g2_dfrbp_1 _12629_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net644),
    .D(net896),
    .Q_N(_05875_),
    .Q(\xdi[7] ));
 sg13g2_dfrbp_1 _12630_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net643),
    .D(_01146_),
    .Q_N(_05874_),
    .Q(\xdi[8] ));
 sg13g2_dfrbp_1 _12631_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net642),
    .D(net917),
    .Q_N(_05873_),
    .Q(\xdi[9] ));
 sg13g2_dfrbp_1 _12632_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net641),
    .D(net907),
    .Q_N(_05872_),
    .Q(\xdi[10] ));
 sg13g2_dfrbp_1 _12633_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net640),
    .D(_01149_),
    .Q_N(_05871_),
    .Q(\xdi[11] ));
 sg13g2_dfrbp_1 _12634_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net639),
    .D(_01150_),
    .Q_N(_05870_),
    .Q(\xdi[12] ));
 sg13g2_dfrbp_1 _12635_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net638),
    .D(net892),
    .Q_N(_05869_),
    .Q(\xdi[13] ));
 sg13g2_dfrbp_1 _12636_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net637),
    .D(_01152_),
    .Q_N(_05868_),
    .Q(\xdi[14] ));
 sg13g2_dfrbp_1 _12637_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net481),
    .D(net920),
    .Q_N(_06034_),
    .Q(\xdi[15] ));
 sg13g2_dfrbp_1 _12638_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net3717),
    .D(_00000_),
    .Q_N(_00544_),
    .Q(\ckd[0] ));
 sg13g2_dfrbp_1 _12639_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net3717),
    .D(_00001_),
    .Q_N(_06035_),
    .Q(\ckd[1] ));
 sg13g2_dfrbp_1 _12640_ (.CLK(clknet_2_2__leaf_jclk_regs),
    .RESET_B(net3717),
    .D(net928),
    .Q_N(_00545_),
    .Q(\ckd[2] ));
 sg13g2_dfrbp_1 _12641_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net543),
    .D(\bsq[1] ),
    .Q_N(_06036_),
    .Q(bsq1r));
 sg13g2_dfrbp_1 _12642_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net3953),
    .D(_00003_),
    .Q_N(_05867_),
    .Q(exintest));
 sg13g2_dfrbp_1 _12643_ (.CLK(net3842),
    .RESET_B(net636),
    .D(_01154_),
    .Q_N(_00221_),
    .Q(\cpu.regs[8][0] ));
 sg13g2_dfrbp_1 _12644_ (.CLK(net3844),
    .RESET_B(net635),
    .D(_01155_),
    .Q_N(_00220_),
    .Q(\cpu.regs[8][1] ));
 sg13g2_dfrbp_1 _12645_ (.CLK(net3795),
    .RESET_B(net634),
    .D(_01156_),
    .Q_N(_00219_),
    .Q(\cpu.regs[8][2] ));
 sg13g2_dfrbp_1 _12646_ (.CLK(net3861),
    .RESET_B(net633),
    .D(_01157_),
    .Q_N(_00218_),
    .Q(\cpu.regs[8][3] ));
 sg13g2_dfrbp_1 _12647_ (.CLK(net3844),
    .RESET_B(net632),
    .D(_01158_),
    .Q_N(_00217_),
    .Q(\cpu.regs[8][4] ));
 sg13g2_dfrbp_1 _12648_ (.CLK(net3868),
    .RESET_B(net631),
    .D(_01159_),
    .Q_N(_00216_),
    .Q(\cpu.regs[8][5] ));
 sg13g2_dfrbp_1 _12649_ (.CLK(net3847),
    .RESET_B(net630),
    .D(_01160_),
    .Q_N(_00215_),
    .Q(\cpu.regs[8][6] ));
 sg13g2_dfrbp_1 _12650_ (.CLK(net3864),
    .RESET_B(net629),
    .D(_01161_),
    .Q_N(_00214_),
    .Q(\cpu.regs[8][7] ));
 sg13g2_dfrbp_1 _12651_ (.CLK(net3867),
    .RESET_B(net628),
    .D(_01162_),
    .Q_N(_00213_),
    .Q(\cpu.regs[8][8] ));
 sg13g2_dfrbp_1 _12652_ (.CLK(net3845),
    .RESET_B(net627),
    .D(_01163_),
    .Q_N(_00212_),
    .Q(\cpu.regs[8][9] ));
 sg13g2_dfrbp_1 _12653_ (.CLK(net3868),
    .RESET_B(net626),
    .D(_01164_),
    .Q_N(_00211_),
    .Q(\cpu.regs[8][10] ));
 sg13g2_dfrbp_1 _12654_ (.CLK(net3857),
    .RESET_B(net625),
    .D(_01165_),
    .Q_N(_00210_),
    .Q(\cpu.regs[8][11] ));
 sg13g2_dfrbp_1 _12655_ (.CLK(net3807),
    .RESET_B(net624),
    .D(_01166_),
    .Q_N(_00209_),
    .Q(\cpu.regs[8][12] ));
 sg13g2_dfrbp_1 _12656_ (.CLK(net3807),
    .RESET_B(net623),
    .D(_01167_),
    .Q_N(_00208_),
    .Q(\cpu.regs[8][13] ));
 sg13g2_dfrbp_1 _12657_ (.CLK(net3854),
    .RESET_B(net622),
    .D(_01168_),
    .Q_N(_00207_),
    .Q(\cpu.regs[8][14] ));
 sg13g2_dfrbp_1 _12658_ (.CLK(net3851),
    .RESET_B(net621),
    .D(_01169_),
    .Q_N(_00206_),
    .Q(\cpu.regs[8][15] ));
 sg13g2_dfrbp_1 _12659_ (.CLK(net3837),
    .RESET_B(net620),
    .D(_01170_),
    .Q_N(_00205_),
    .Q(\cpu.regs[8][16] ));
 sg13g2_dfrbp_1 _12660_ (.CLK(net3859),
    .RESET_B(net619),
    .D(_01171_),
    .Q_N(_00204_),
    .Q(\cpu.regs[8][17] ));
 sg13g2_dfrbp_1 _12661_ (.CLK(net3832),
    .RESET_B(net618),
    .D(_01172_),
    .Q_N(_00203_),
    .Q(\cpu.regs[8][18] ));
 sg13g2_dfrbp_1 _12662_ (.CLK(net3830),
    .RESET_B(net617),
    .D(_01173_),
    .Q_N(_00202_),
    .Q(\cpu.regs[8][19] ));
 sg13g2_dfrbp_1 _12663_ (.CLK(net3803),
    .RESET_B(net616),
    .D(_01174_),
    .Q_N(_00201_),
    .Q(\cpu.regs[8][20] ));
 sg13g2_dfrbp_1 _12664_ (.CLK(net3819),
    .RESET_B(net615),
    .D(_01175_),
    .Q_N(_00200_),
    .Q(\cpu.regs[8][21] ));
 sg13g2_dfrbp_1 _12665_ (.CLK(net3814),
    .RESET_B(net614),
    .D(_01176_),
    .Q_N(_00199_),
    .Q(\cpu.regs[8][22] ));
 sg13g2_dfrbp_1 _12666_ (.CLK(net3814),
    .RESET_B(net613),
    .D(_01177_),
    .Q_N(_00198_),
    .Q(\cpu.regs[8][23] ));
 sg13g2_dfrbp_1 _12667_ (.CLK(net3813),
    .RESET_B(net612),
    .D(_01178_),
    .Q_N(_00197_),
    .Q(\cpu.regs[8][24] ));
 sg13g2_dfrbp_1 _12668_ (.CLK(net3821),
    .RESET_B(net611),
    .D(_01179_),
    .Q_N(_00196_),
    .Q(\cpu.regs[8][25] ));
 sg13g2_dfrbp_1 _12669_ (.CLK(net3804),
    .RESET_B(net610),
    .D(_01180_),
    .Q_N(_00195_),
    .Q(\cpu.regs[8][26] ));
 sg13g2_dfrbp_1 _12670_ (.CLK(net3817),
    .RESET_B(net609),
    .D(_01181_),
    .Q_N(_00194_),
    .Q(\cpu.regs[8][27] ));
 sg13g2_dfrbp_1 _12671_ (.CLK(net3824),
    .RESET_B(net608),
    .D(_01182_),
    .Q_N(_00193_),
    .Q(\cpu.regs[8][28] ));
 sg13g2_dfrbp_1 _12672_ (.CLK(net3826),
    .RESET_B(net607),
    .D(_01183_),
    .Q_N(_00192_),
    .Q(\cpu.regs[8][29] ));
 sg13g2_dfrbp_1 _12673_ (.CLK(net3807),
    .RESET_B(net606),
    .D(_01184_),
    .Q_N(_00191_),
    .Q(\cpu.regs[8][30] ));
 sg13g2_dfrbp_1 _12674_ (.CLK(net3802),
    .RESET_B(net605),
    .D(_01185_),
    .Q_N(_00190_),
    .Q(\cpu.regs[8][31] ));
 sg13g2_dfrbp_1 _12675_ (.CLK(net3840),
    .RESET_B(net604),
    .D(_01186_),
    .Q_N(_00189_),
    .Q(\cpu.regs[15][0] ));
 sg13g2_dfrbp_1 _12676_ (.CLK(net3841),
    .RESET_B(net603),
    .D(_01187_),
    .Q_N(_00188_),
    .Q(\cpu.regs[15][1] ));
 sg13g2_dfrbp_1 _12677_ (.CLK(net3840),
    .RESET_B(net602),
    .D(_01188_),
    .Q_N(_00187_),
    .Q(\cpu.regs[15][2] ));
 sg13g2_dfrbp_1 _12678_ (.CLK(net3854),
    .RESET_B(net601),
    .D(_01189_),
    .Q_N(_00186_),
    .Q(\cpu.regs[15][3] ));
 sg13g2_dfrbp_1 _12679_ (.CLK(net3840),
    .RESET_B(net600),
    .D(_01190_),
    .Q_N(_00185_),
    .Q(\cpu.regs[15][4] ));
 sg13g2_dfrbp_1 _12680_ (.CLK(net3868),
    .RESET_B(net599),
    .D(_01191_),
    .Q_N(_00184_),
    .Q(\cpu.regs[15][5] ));
 sg13g2_dfrbp_1 _12681_ (.CLK(net3847),
    .RESET_B(net598),
    .D(_01192_),
    .Q_N(_00183_),
    .Q(\cpu.regs[15][6] ));
 sg13g2_dfrbp_1 _12682_ (.CLK(net3862),
    .RESET_B(net597),
    .D(_01193_),
    .Q_N(_00182_),
    .Q(\cpu.regs[15][7] ));
 sg13g2_dfrbp_1 _12683_ (.CLK(net3866),
    .RESET_B(net596),
    .D(_01194_),
    .Q_N(_00181_),
    .Q(\cpu.regs[15][8] ));
 sg13g2_dfrbp_1 _12684_ (.CLK(net3845),
    .RESET_B(net595),
    .D(_01195_),
    .Q_N(_00180_),
    .Q(\cpu.regs[15][9] ));
 sg13g2_dfrbp_1 _12685_ (.CLK(net3867),
    .RESET_B(net594),
    .D(_01196_),
    .Q_N(_00179_),
    .Q(\cpu.regs[15][10] ));
 sg13g2_dfrbp_1 _12686_ (.CLK(net3856),
    .RESET_B(net593),
    .D(_01197_),
    .Q_N(_00178_),
    .Q(\cpu.regs[15][11] ));
 sg13g2_dfrbp_1 _12687_ (.CLK(net3807),
    .RESET_B(net592),
    .D(_01198_),
    .Q_N(_00177_),
    .Q(\cpu.regs[15][12] ));
 sg13g2_dfrbp_1 _12688_ (.CLK(net3806),
    .RESET_B(net591),
    .D(_01199_),
    .Q_N(_00176_),
    .Q(\cpu.regs[15][13] ));
 sg13g2_dfrbp_1 _12689_ (.CLK(net3854),
    .RESET_B(net590),
    .D(_01200_),
    .Q_N(_00175_),
    .Q(\cpu.regs[15][14] ));
 sg13g2_dfrbp_1 _12690_ (.CLK(net3852),
    .RESET_B(net589),
    .D(_01201_),
    .Q_N(_00174_),
    .Q(\cpu.regs[15][15] ));
 sg13g2_dfrbp_1 _12691_ (.CLK(net3834),
    .RESET_B(net588),
    .D(_01202_),
    .Q_N(_00173_),
    .Q(\cpu.regs[15][16] ));
 sg13g2_dfrbp_1 _12692_ (.CLK(net3858),
    .RESET_B(net587),
    .D(_01203_),
    .Q_N(_00172_),
    .Q(\cpu.regs[15][17] ));
 sg13g2_dfrbp_1 _12693_ (.CLK(net3829),
    .RESET_B(net586),
    .D(_01204_),
    .Q_N(_00171_),
    .Q(\cpu.regs[15][18] ));
 sg13g2_dfrbp_1 _12694_ (.CLK(net3830),
    .RESET_B(net585),
    .D(_01205_),
    .Q_N(_00170_),
    .Q(\cpu.regs[15][19] ));
 sg13g2_dfrbp_1 _12695_ (.CLK(net3803),
    .RESET_B(net584),
    .D(_01206_),
    .Q_N(_00169_),
    .Q(\cpu.regs[15][20] ));
 sg13g2_dfrbp_1 _12696_ (.CLK(net3821),
    .RESET_B(net583),
    .D(_01207_),
    .Q_N(_00168_),
    .Q(\cpu.regs[15][21] ));
 sg13g2_dfrbp_1 _12697_ (.CLK(net3814),
    .RESET_B(net582),
    .D(_01208_),
    .Q_N(_00167_),
    .Q(\cpu.regs[15][22] ));
 sg13g2_dfrbp_1 _12698_ (.CLK(net3820),
    .RESET_B(net581),
    .D(_01209_),
    .Q_N(_00166_),
    .Q(\cpu.regs[15][23] ));
 sg13g2_dfrbp_1 _12699_ (.CLK(net3816),
    .RESET_B(net580),
    .D(_01210_),
    .Q_N(_00165_),
    .Q(\cpu.regs[15][24] ));
 sg13g2_dfrbp_1 _12700_ (.CLK(net3832),
    .RESET_B(net579),
    .D(_01211_),
    .Q_N(_00164_),
    .Q(\cpu.regs[15][25] ));
 sg13g2_dfrbp_1 _12701_ (.CLK(net3813),
    .RESET_B(net578),
    .D(_01212_),
    .Q_N(_00163_),
    .Q(\cpu.regs[15][26] ));
 sg13g2_dfrbp_1 _12702_ (.CLK(net3825),
    .RESET_B(net577),
    .D(_01213_),
    .Q_N(_00162_),
    .Q(\cpu.regs[15][27] ));
 sg13g2_dfrbp_1 _12703_ (.CLK(net3817),
    .RESET_B(net576),
    .D(_01214_),
    .Q_N(_00161_),
    .Q(\cpu.regs[15][28] ));
 sg13g2_dfrbp_1 _12704_ (.CLK(net3827),
    .RESET_B(net575),
    .D(_01215_),
    .Q_N(_00160_),
    .Q(\cpu.regs[15][29] ));
 sg13g2_dfrbp_1 _12705_ (.CLK(net3810),
    .RESET_B(net574),
    .D(_01216_),
    .Q_N(_00159_),
    .Q(\cpu.regs[15][30] ));
 sg13g2_dfrbp_1 _12706_ (.CLK(net3813),
    .RESET_B(net573),
    .D(_01217_),
    .Q_N(_00158_),
    .Q(\cpu.regs[15][31] ));
 sg13g2_dfrbp_1 _12707_ (.CLK(net3842),
    .RESET_B(net572),
    .D(_01218_),
    .Q_N(_00157_),
    .Q(\cpu.regs[9][0] ));
 sg13g2_dfrbp_1 _12708_ (.CLK(net3841),
    .RESET_B(net571),
    .D(_01219_),
    .Q_N(_00156_),
    .Q(\cpu.regs[9][1] ));
 sg13g2_dfrbp_1 _12709_ (.CLK(net3795),
    .RESET_B(net570),
    .D(_01220_),
    .Q_N(_00155_),
    .Q(\cpu.regs[9][2] ));
 sg13g2_dfrbp_1 _12710_ (.CLK(net3862),
    .RESET_B(net569),
    .D(_01221_),
    .Q_N(_00154_),
    .Q(\cpu.regs[9][3] ));
 sg13g2_dfrbp_1 _12711_ (.CLK(net3796),
    .RESET_B(net568),
    .D(_01222_),
    .Q_N(_00153_),
    .Q(\cpu.regs[9][4] ));
 sg13g2_dfrbp_1 _12712_ (.CLK(net3868),
    .RESET_B(net567),
    .D(_01223_),
    .Q_N(_00152_),
    .Q(\cpu.regs[9][5] ));
 sg13g2_dfrbp_1 _12713_ (.CLK(net3847),
    .RESET_B(net566),
    .D(_01224_),
    .Q_N(_00151_),
    .Q(\cpu.regs[9][6] ));
 sg13g2_dfrbp_1 _12714_ (.CLK(net3865),
    .RESET_B(net565),
    .D(_01225_),
    .Q_N(_00150_),
    .Q(\cpu.regs[9][7] ));
 sg13g2_dfrbp_1 _12715_ (.CLK(net3867),
    .RESET_B(net564),
    .D(_01226_),
    .Q_N(_00149_),
    .Q(\cpu.regs[9][8] ));
 sg13g2_dfrbp_1 _12716_ (.CLK(net3845),
    .RESET_B(net563),
    .D(_01227_),
    .Q_N(_00148_),
    .Q(\cpu.regs[9][9] ));
 sg13g2_dfrbp_1 _12717_ (.CLK(net3858),
    .RESET_B(net562),
    .D(_01228_),
    .Q_N(_00147_),
    .Q(\cpu.regs[9][10] ));
 sg13g2_dfrbp_1 _12718_ (.CLK(net3856),
    .RESET_B(net561),
    .D(_01229_),
    .Q_N(_00146_),
    .Q(\cpu.regs[9][11] ));
 sg13g2_dfrbp_1 _12719_ (.CLK(net3804),
    .RESET_B(net560),
    .D(_01230_),
    .Q_N(_00145_),
    .Q(\cpu.regs[9][12] ));
 sg13g2_dfrbp_1 _12720_ (.CLK(net3806),
    .RESET_B(net559),
    .D(_01231_),
    .Q_N(_00144_),
    .Q(\cpu.regs[9][13] ));
 sg13g2_dfrbp_1 _12721_ (.CLK(net3854),
    .RESET_B(net558),
    .D(_01232_),
    .Q_N(_00143_),
    .Q(\cpu.regs[9][14] ));
 sg13g2_dfrbp_1 _12722_ (.CLK(net3851),
    .RESET_B(net557),
    .D(_01233_),
    .Q_N(_00142_),
    .Q(\cpu.regs[9][15] ));
 sg13g2_dfrbp_1 _12723_ (.CLK(net3837),
    .RESET_B(net556),
    .D(_01234_),
    .Q_N(_00141_),
    .Q(\cpu.regs[9][16] ));
 sg13g2_dfrbp_1 _12724_ (.CLK(net3859),
    .RESET_B(net555),
    .D(_01235_),
    .Q_N(_00140_),
    .Q(\cpu.regs[9][17] ));
 sg13g2_dfrbp_1 _12725_ (.CLK(net3831),
    .RESET_B(net554),
    .D(_01236_),
    .Q_N(_00139_),
    .Q(\cpu.regs[9][18] ));
 sg13g2_dfrbp_1 _12726_ (.CLK(net3830),
    .RESET_B(net553),
    .D(_01237_),
    .Q_N(_00138_),
    .Q(\cpu.regs[9][19] ));
 sg13g2_dfrbp_1 _12727_ (.CLK(net3803),
    .RESET_B(net552),
    .D(_01238_),
    .Q_N(_00137_),
    .Q(\cpu.regs[9][20] ));
 sg13g2_dfrbp_1 _12728_ (.CLK(net3819),
    .RESET_B(net551),
    .D(_01239_),
    .Q_N(_00136_),
    .Q(\cpu.regs[9][21] ));
 sg13g2_dfrbp_1 _12729_ (.CLK(net3814),
    .RESET_B(net550),
    .D(_01240_),
    .Q_N(_00135_),
    .Q(\cpu.regs[9][22] ));
 sg13g2_dfrbp_1 _12730_ (.CLK(net3818),
    .RESET_B(net549),
    .D(_01241_),
    .Q_N(_00134_),
    .Q(\cpu.regs[9][23] ));
 sg13g2_dfrbp_1 _12731_ (.CLK(net3813),
    .RESET_B(net548),
    .D(_01242_),
    .Q_N(_00133_),
    .Q(\cpu.regs[9][24] ));
 sg13g2_dfrbp_1 _12732_ (.CLK(net3829),
    .RESET_B(net547),
    .D(_01243_),
    .Q_N(_00132_),
    .Q(\cpu.regs[9][25] ));
 sg13g2_dfrbp_1 _12733_ (.CLK(net3804),
    .RESET_B(net546),
    .D(_01244_),
    .Q_N(_00131_),
    .Q(\cpu.regs[9][26] ));
 sg13g2_dfrbp_1 _12734_ (.CLK(net3817),
    .RESET_B(net545),
    .D(_01245_),
    .Q_N(_00130_),
    .Q(\cpu.regs[9][27] ));
 sg13g2_dfrbp_1 _12735_ (.CLK(net3824),
    .RESET_B(net544),
    .D(_01246_),
    .Q_N(_00129_),
    .Q(\cpu.regs[9][28] ));
 sg13g2_dfrbp_1 _12736_ (.CLK(net3826),
    .RESET_B(net542),
    .D(_01247_),
    .Q_N(_00128_),
    .Q(\cpu.regs[9][29] ));
 sg13g2_dfrbp_1 _12737_ (.CLK(net3809),
    .RESET_B(net541),
    .D(_01248_),
    .Q_N(_00127_),
    .Q(\cpu.regs[9][30] ));
 sg13g2_dfrbp_1 _12738_ (.CLK(net3802),
    .RESET_B(net540),
    .D(_01249_),
    .Q_N(_00126_),
    .Q(\cpu.regs[9][31] ));
 sg13g2_dfrbp_1 _12739_ (.CLK(_00591_),
    .RESET_B(net1),
    .D(_01535_),
    .Q_N(_05866_),
    .Q(\jtag0.tapst[0] ));
 sg13g2_dfrbp_1 _12740_ (.CLK(_00592_),
    .RESET_B(net1),
    .D(_01536_),
    .Q_N(_05865_),
    .Q(\jtag0.tapst[1] ));
 sg13g2_dfrbp_1 _12741_ (.CLK(_00593_),
    .RESET_B(net3953),
    .D(_01537_),
    .Q_N(_05864_),
    .Q(\jtag0.tapst[2] ));
 sg13g2_dfrbp_1 _12742_ (.CLK(_00594_),
    .RESET_B(net3953),
    .D(_01538_),
    .Q_N(_06037_),
    .Q(\jtag0.tapst[3] ));
 sg13g2_dfrbp_1 _12743_ (.CLK(net3941),
    .RESET_B(net539),
    .D(net3),
    .Q_N(_05863_),
    .Q(\jtag0.stdi ));
 sg13g2_dfrbp_1 _12744_ (.CLK(_00595_),
    .RESET_B(net3953),
    .D(_01250_),
    .Q_N(_05862_),
    .Q(\jtag0.ir[0] ));
 sg13g2_dfrbp_1 _12745_ (.CLK(_00596_),
    .RESET_B(net3953),
    .D(_01251_),
    .Q_N(_05861_),
    .Q(\jtag0.ir[1] ));
 sg13g2_dfrbp_1 _12746_ (.CLK(_00597_),
    .RESET_B(net3953),
    .D(_01252_),
    .Q_N(_00125_),
    .Q(\jtag0.ir[2] ));
 sg13g2_dfrbp_1 _12747_ (.CLK(_00598_),
    .RESET_B(net727),
    .D(_01253_),
    .Q_N(_06038_),
    .Q(\jtag0.byp ));
 sg13g2_dfrbp_1 _12748_ (.CLK(net3941),
    .RESET_B(net535),
    .D(net2),
    .Q_N(_00124_),
    .Q(\jtag0.stms ));
 sg13g2_dfrbp_1 _12749_ (.CLK(_00599_),
    .RESET_B(net533),
    .D(_01254_),
    .Q_N(_05860_),
    .Q(\jtag0.idr[0] ));
 sg13g2_dfrbp_1 _12750_ (.CLK(_00600_),
    .RESET_B(net530),
    .D(_01255_),
    .Q_N(_05859_),
    .Q(\jtag0.idr[1] ));
 sg13g2_dfrbp_1 _12751_ (.CLK(_00601_),
    .RESET_B(net527),
    .D(_01256_),
    .Q_N(_05858_),
    .Q(\jtag0.idr[2] ));
 sg13g2_dfrbp_1 _12752_ (.CLK(_00602_),
    .RESET_B(net524),
    .D(_01257_),
    .Q_N(_05857_),
    .Q(\jtag0.idr[3] ));
 sg13g2_dfrbp_1 _12753_ (.CLK(_00603_),
    .RESET_B(net521),
    .D(_01258_),
    .Q_N(_05856_),
    .Q(\jtag0.idr[4] ));
 sg13g2_dfrbp_1 _12754_ (.CLK(_00604_),
    .RESET_B(net518),
    .D(_01259_),
    .Q_N(_05855_),
    .Q(\jtag0.idr[5] ));
 sg13g2_dfrbp_1 _12755_ (.CLK(_00605_),
    .RESET_B(net515),
    .D(_01260_),
    .Q_N(_05854_),
    .Q(\jtag0.idr[6] ));
 sg13g2_dfrbp_1 _12756_ (.CLK(_00606_),
    .RESET_B(net513),
    .D(_01261_),
    .Q_N(_05853_),
    .Q(\jtag0.idr[7] ));
 sg13g2_dfrbp_1 _12757_ (.CLK(_00607_),
    .RESET_B(net512),
    .D(_01262_),
    .Q_N(_05852_),
    .Q(\jtag0.idr[8] ));
 sg13g2_dfrbp_1 _12758_ (.CLK(_00608_),
    .RESET_B(net509),
    .D(_01263_),
    .Q_N(_05851_),
    .Q(\jtag0.idr[9] ));
 sg13g2_dfrbp_1 _12759_ (.CLK(_00609_),
    .RESET_B(net506),
    .D(_01264_),
    .Q_N(_05850_),
    .Q(\jtag0.idr[10] ));
 sg13g2_dfrbp_1 _12760_ (.CLK(_00610_),
    .RESET_B(net503),
    .D(_01265_),
    .Q_N(_05849_),
    .Q(\jtag0.idr[11] ));
 sg13g2_dfrbp_1 _12761_ (.CLK(_00611_),
    .RESET_B(net500),
    .D(_01266_),
    .Q_N(_05848_),
    .Q(\jtag0.idr[12] ));
 sg13g2_dfrbp_1 _12762_ (.CLK(_00612_),
    .RESET_B(net499),
    .D(_01267_),
    .Q_N(_05847_),
    .Q(\jtag0.idr[13] ));
 sg13g2_dfrbp_1 _12763_ (.CLK(_00613_),
    .RESET_B(net498),
    .D(_01268_),
    .Q_N(_05846_),
    .Q(\jtag0.idr[14] ));
 sg13g2_dfrbp_1 _12764_ (.CLK(_00614_),
    .RESET_B(net497),
    .D(_01269_),
    .Q_N(_05845_),
    .Q(\jtag0.idr[15] ));
 sg13g2_dfrbp_1 _12765_ (.CLK(_00615_),
    .RESET_B(net496),
    .D(_01270_),
    .Q_N(_05844_),
    .Q(\jtag0.idr[16] ));
 sg13g2_dfrbp_1 _12766_ (.CLK(_00616_),
    .RESET_B(net495),
    .D(_01271_),
    .Q_N(_05843_),
    .Q(\jtag0.idr[17] ));
 sg13g2_dfrbp_1 _12767_ (.CLK(_00617_),
    .RESET_B(net494),
    .D(_01272_),
    .Q_N(_05842_),
    .Q(\jtag0.idr[18] ));
 sg13g2_dfrbp_1 _12768_ (.CLK(_00618_),
    .RESET_B(net493),
    .D(_01273_),
    .Q_N(_05841_),
    .Q(\jtag0.idr[19] ));
 sg13g2_dfrbp_1 _12769_ (.CLK(_00619_),
    .RESET_B(net492),
    .D(_01274_),
    .Q_N(_05840_),
    .Q(\jtag0.idr[20] ));
 sg13g2_dfrbp_1 _12770_ (.CLK(_00620_),
    .RESET_B(net491),
    .D(_01275_),
    .Q_N(_05839_),
    .Q(\jtag0.idr[21] ));
 sg13g2_dfrbp_1 _12771_ (.CLK(_00621_),
    .RESET_B(net490),
    .D(_01276_),
    .Q_N(_05838_),
    .Q(\jtag0.idr[22] ));
 sg13g2_dfrbp_1 _12772_ (.CLK(_00622_),
    .RESET_B(net489),
    .D(_01277_),
    .Q_N(_05837_),
    .Q(\jtag0.idr[23] ));
 sg13g2_dfrbp_1 _12773_ (.CLK(_00623_),
    .RESET_B(net488),
    .D(_01278_),
    .Q_N(_05836_),
    .Q(\jtag0.idr[24] ));
 sg13g2_dfrbp_1 _12774_ (.CLK(_00624_),
    .RESET_B(net487),
    .D(_01279_),
    .Q_N(_05835_),
    .Q(\jtag0.idr[25] ));
 sg13g2_dfrbp_1 _12775_ (.CLK(_00625_),
    .RESET_B(net486),
    .D(_01280_),
    .Q_N(_05834_),
    .Q(\jtag0.idr[26] ));
 sg13g2_dfrbp_1 _12776_ (.CLK(_00626_),
    .RESET_B(net485),
    .D(_01281_),
    .Q_N(_05833_),
    .Q(\jtag0.idr[27] ));
 sg13g2_dfrbp_1 _12777_ (.CLK(_00627_),
    .RESET_B(net482),
    .D(_01282_),
    .Q_N(_05832_),
    .Q(\jtag0.idr[28] ));
 sg13g2_dfrbp_1 _12778_ (.CLK(_00628_),
    .RESET_B(net478),
    .D(_01283_),
    .Q_N(_05831_),
    .Q(\jtag0.idr[29] ));
 sg13g2_dfrbp_1 _12779_ (.CLK(_00629_),
    .RESET_B(net475),
    .D(_01284_),
    .Q_N(_05830_),
    .Q(\jtag0.idr[30] ));
 sg13g2_dfrbp_1 _12780_ (.CLK(_00630_),
    .RESET_B(net472),
    .D(_01285_),
    .Q_N(_05829_),
    .Q(\jtag0.idr[31] ));
 sg13g2_dfrbp_1 _12781_ (.CLK(_00631_),
    .RESET_B(net469),
    .D(_01286_),
    .Q_N(_05828_),
    .Q(\jtag0.bssh[0] ));
 sg13g2_dfrbp_1 _12782_ (.CLK(_00632_),
    .RESET_B(net467),
    .D(_01287_),
    .Q_N(_05827_),
    .Q(\jtag0.bssh[1] ));
 sg13g2_dfrbp_1 _12783_ (.CLK(_00633_),
    .RESET_B(net465),
    .D(_01288_),
    .Q_N(_05826_),
    .Q(\jtag0.bssh[2] ));
 sg13g2_dfrbp_1 _12784_ (.CLK(_00634_),
    .RESET_B(net463),
    .D(_01289_),
    .Q_N(_05825_),
    .Q(\jtag0.bssh[3] ));
 sg13g2_dfrbp_1 _12785_ (.CLK(_00635_),
    .RESET_B(net461),
    .D(_01290_),
    .Q_N(_05824_),
    .Q(\jtag0.bssh[4] ));
 sg13g2_dfrbp_1 _12786_ (.CLK(_00636_),
    .RESET_B(net459),
    .D(_01291_),
    .Q_N(_05823_),
    .Q(\jtag0.bssh[5] ));
 sg13g2_dfrbp_1 _12787_ (.CLK(_00637_),
    .RESET_B(net457),
    .D(_01292_),
    .Q_N(_05822_),
    .Q(\jtag0.bssh[6] ));
 sg13g2_dfrbp_1 _12788_ (.CLK(_00638_),
    .RESET_B(net455),
    .D(_01293_),
    .Q_N(_05821_),
    .Q(\jtag0.bssh[7] ));
 sg13g2_dfrbp_1 _12789_ (.CLK(_00639_),
    .RESET_B(net453),
    .D(_01294_),
    .Q_N(_05820_),
    .Q(\jtag0.bssh[8] ));
 sg13g2_dfrbp_1 _12790_ (.CLK(_00640_),
    .RESET_B(net451),
    .D(_01295_),
    .Q_N(_05819_),
    .Q(\jtag0.bssh[9] ));
 sg13g2_dfrbp_1 _12791_ (.CLK(_00641_),
    .RESET_B(net449),
    .D(_01296_),
    .Q_N(_05818_),
    .Q(\jtag0.bssh[10] ));
 sg13g2_dfrbp_1 _12792_ (.CLK(_00642_),
    .RESET_B(net447),
    .D(_01297_),
    .Q_N(_05817_),
    .Q(\jtag0.bssh[11] ));
 sg13g2_dfrbp_1 _12793_ (.CLK(_00643_),
    .RESET_B(net445),
    .D(_01298_),
    .Q_N(_05816_),
    .Q(\jtag0.bssh[12] ));
 sg13g2_dfrbp_1 _12794_ (.CLK(_00644_),
    .RESET_B(net443),
    .D(_01299_),
    .Q_N(_05815_),
    .Q(\jtag0.bssh[13] ));
 sg13g2_dfrbp_1 _12795_ (.CLK(_00645_),
    .RESET_B(net441),
    .D(_01300_),
    .Q_N(_05814_),
    .Q(\jtag0.bssh[14] ));
 sg13g2_dfrbp_1 _12796_ (.CLK(_00646_),
    .RESET_B(net439),
    .D(_01301_),
    .Q_N(_05813_),
    .Q(\jtag0.bssh[15] ));
 sg13g2_dfrbp_1 _12797_ (.CLK(_00647_),
    .RESET_B(net437),
    .D(_01302_),
    .Q_N(_05812_),
    .Q(\jtag0.bssh[16] ));
 sg13g2_dfrbp_1 _12798_ (.CLK(_00648_),
    .RESET_B(net435),
    .D(_01303_),
    .Q_N(_05811_),
    .Q(\jtag0.bssh[17] ));
 sg13g2_dfrbp_1 _12799_ (.CLK(_00649_),
    .RESET_B(net433),
    .D(_01304_),
    .Q_N(_05810_),
    .Q(\jtag0.bssh[18] ));
 sg13g2_dfrbp_1 _12800_ (.CLK(_00650_),
    .RESET_B(net431),
    .D(_01305_),
    .Q_N(_05809_),
    .Q(\jtag0.bssh[19] ));
 sg13g2_dfrbp_1 _12801_ (.CLK(_00651_),
    .RESET_B(net429),
    .D(_01306_),
    .Q_N(_05808_),
    .Q(\jtag0.bssh[20] ));
 sg13g2_dfrbp_1 _12802_ (.CLK(_00652_),
    .RESET_B(net428),
    .D(_01307_),
    .Q_N(_05807_),
    .Q(\jtag0.bssh[21] ));
 sg13g2_dfrbp_1 _12803_ (.CLK(_00653_),
    .RESET_B(net427),
    .D(_01308_),
    .Q_N(_05806_),
    .Q(\jtag0.bssh[22] ));
 sg13g2_dfrbp_1 _12804_ (.CLK(_00654_),
    .RESET_B(net426),
    .D(_01309_),
    .Q_N(_05805_),
    .Q(\jtag0.bssh[23] ));
 sg13g2_dfrbp_1 _12805_ (.CLK(_00655_),
    .RESET_B(net425),
    .D(_01310_),
    .Q_N(_05804_),
    .Q(\jtag0.bssh[24] ));
 sg13g2_dfrbp_1 _12806_ (.CLK(_00656_),
    .RESET_B(net424),
    .D(_01311_),
    .Q_N(_05803_),
    .Q(\jtag0.bssh[25] ));
 sg13g2_dfrbp_1 _12807_ (.CLK(_00657_),
    .RESET_B(net423),
    .D(_01312_),
    .Q_N(_05802_),
    .Q(\jtag0.bssh[26] ));
 sg13g2_dfrbp_1 _12808_ (.CLK(_00658_),
    .RESET_B(net422),
    .D(_01313_),
    .Q_N(_05801_),
    .Q(\jtag0.bssh[27] ));
 sg13g2_dfrbp_1 _12809_ (.CLK(_00659_),
    .RESET_B(net421),
    .D(_01314_),
    .Q_N(_05800_),
    .Q(\jtag0.bssh[28] ));
 sg13g2_dfrbp_1 _12810_ (.CLK(_00660_),
    .RESET_B(net420),
    .D(_01315_),
    .Q_N(_05799_),
    .Q(\jtag0.bssh[29] ));
 sg13g2_dfrbp_1 _12811_ (.CLK(_00661_),
    .RESET_B(net419),
    .D(_01316_),
    .Q_N(_05798_),
    .Q(\bsq[0] ));
 sg13g2_dfrbp_1 _12812_ (.CLK(_00662_),
    .RESET_B(net417),
    .D(_01317_),
    .Q_N(_05797_),
    .Q(\bsq[1] ));
 sg13g2_dfrbp_1 _12813_ (.CLK(_00663_),
    .RESET_B(net415),
    .D(_01318_),
    .Q_N(_05796_),
    .Q(\bsq[2] ));
 sg13g2_dfrbp_1 _12814_ (.CLK(_00664_),
    .RESET_B(net414),
    .D(_01319_),
    .Q_N(_05795_),
    .Q(\bsq[3] ));
 sg13g2_dfrbp_1 _12815_ (.CLK(_00665_),
    .RESET_B(net413),
    .D(_01320_),
    .Q_N(_05794_),
    .Q(\bsq[4] ));
 sg13g2_dfrbp_1 _12816_ (.CLK(_00666_),
    .RESET_B(net411),
    .D(_01321_),
    .Q_N(_05793_),
    .Q(\bsq[5] ));
 sg13g2_dfrbp_1 _12817_ (.CLK(_00667_),
    .RESET_B(net409),
    .D(_01322_),
    .Q_N(_05792_),
    .Q(\bsq[6] ));
 sg13g2_dfrbp_1 _12818_ (.CLK(_00668_),
    .RESET_B(net408),
    .D(_01323_),
    .Q_N(_05791_),
    .Q(\bsq[7] ));
 sg13g2_dfrbp_1 _12819_ (.CLK(_00669_),
    .RESET_B(net406),
    .D(_01324_),
    .Q_N(_05790_),
    .Q(\bsq[8] ));
 sg13g2_dfrbp_1 _12820_ (.CLK(_00670_),
    .RESET_B(net405),
    .D(_01325_),
    .Q_N(_05789_),
    .Q(\bsq[9] ));
 sg13g2_dfrbp_1 _12821_ (.CLK(_00671_),
    .RESET_B(net403),
    .D(_01326_),
    .Q_N(_05788_),
    .Q(\bsq[10] ));
 sg13g2_dfrbp_1 _12822_ (.CLK(_00672_),
    .RESET_B(net402),
    .D(_01327_),
    .Q_N(_05787_),
    .Q(\bsq[11] ));
 sg13g2_dfrbp_1 _12823_ (.CLK(_00673_),
    .RESET_B(net400),
    .D(_01328_),
    .Q_N(_05786_),
    .Q(\bsq[12] ));
 sg13g2_dfrbp_1 _12824_ (.CLK(_00674_),
    .RESET_B(net398),
    .D(_01329_),
    .Q_N(_05785_),
    .Q(\bsq[13] ));
 sg13g2_dfrbp_1 _12825_ (.CLK(_00675_),
    .RESET_B(net397),
    .D(_01330_),
    .Q_N(_05784_),
    .Q(\bsq[14] ));
 sg13g2_dfrbp_1 _12826_ (.CLK(_00676_),
    .RESET_B(net396),
    .D(_01331_),
    .Q_N(_05783_),
    .Q(\bsq[15] ));
 sg13g2_dfrbp_1 _12827_ (.CLK(_00677_),
    .RESET_B(net394),
    .D(_01332_),
    .Q_N(_05782_),
    .Q(\bsq[16] ));
 sg13g2_dfrbp_1 _12828_ (.CLK(_00678_),
    .RESET_B(net392),
    .D(_01333_),
    .Q_N(_05781_),
    .Q(\bsq[17] ));
 sg13g2_dfrbp_1 _12829_ (.CLK(_00679_),
    .RESET_B(net390),
    .D(_01334_),
    .Q_N(_05780_),
    .Q(\bsq[18] ));
 sg13g2_dfrbp_1 _12830_ (.CLK(_00680_),
    .RESET_B(net389),
    .D(_01335_),
    .Q_N(_05779_),
    .Q(\bsq[19] ));
 sg13g2_dfrbp_1 _12831_ (.CLK(_00681_),
    .RESET_B(net388),
    .D(_01336_),
    .Q_N(_05778_),
    .Q(\bsq[20] ));
 sg13g2_dfrbp_1 _12832_ (.CLK(_00682_),
    .RESET_B(net386),
    .D(_01337_),
    .Q_N(_05777_),
    .Q(\bsq[21] ));
 sg13g2_dfrbp_1 _12833_ (.CLK(_00683_),
    .RESET_B(net385),
    .D(_01338_),
    .Q_N(_05776_),
    .Q(\bsq[22] ));
 sg13g2_dfrbp_1 _12834_ (.CLK(_00684_),
    .RESET_B(net384),
    .D(_01339_),
    .Q_N(_05775_),
    .Q(\bsq[23] ));
 sg13g2_dfrbp_1 _12835_ (.CLK(_00685_),
    .RESET_B(net382),
    .D(_01340_),
    .Q_N(_05774_),
    .Q(\bsq[24] ));
 sg13g2_dfrbp_1 _12836_ (.CLK(_00686_),
    .RESET_B(net381),
    .D(_01341_),
    .Q_N(_05773_),
    .Q(\bsq[25] ));
 sg13g2_dfrbp_1 _12837_ (.CLK(_00687_),
    .RESET_B(net380),
    .D(_01342_),
    .Q_N(_05772_),
    .Q(\bsq[26] ));
 sg13g2_dfrbp_1 _12838_ (.CLK(_00688_),
    .RESET_B(net379),
    .D(_01343_),
    .Q_N(_05771_),
    .Q(\bsq[27] ));
 sg13g2_dfrbp_1 _12839_ (.CLK(_00689_),
    .RESET_B(net378),
    .D(_01344_),
    .Q_N(_05770_),
    .Q(\bsq[28] ));
 sg13g2_dfrbp_1 _12840_ (.CLK(_00690_),
    .RESET_B(net377),
    .D(_01345_),
    .Q_N(_05769_),
    .Q(\bsq[29] ));
 sg13g2_dfrbp_1 _12841_ (.CLK(net3792),
    .RESET_B(net376),
    .D(_01346_),
    .Q_N(_05768_),
    .Q(\cpu.PCreg1[2] ));
 sg13g2_dfrbp_1 _12842_ (.CLK(net3787),
    .RESET_B(net375),
    .D(_01347_),
    .Q_N(_05767_),
    .Q(\cpu.PCreg1[3] ));
 sg13g2_dfrbp_1 _12843_ (.CLK(net3786),
    .RESET_B(net374),
    .D(_01348_),
    .Q_N(_05766_),
    .Q(\cpu.PCreg1[4] ));
 sg13g2_dfrbp_1 _12844_ (.CLK(net3787),
    .RESET_B(net373),
    .D(_01349_),
    .Q_N(_05765_),
    .Q(\cpu.PCreg1[5] ));
 sg13g2_dfrbp_1 _12845_ (.CLK(net3781),
    .RESET_B(net372),
    .D(_01350_),
    .Q_N(_05764_),
    .Q(\cpu.PCreg1[6] ));
 sg13g2_dfrbp_1 _12846_ (.CLK(net3759),
    .RESET_B(net371),
    .D(_01351_),
    .Q_N(_05763_),
    .Q(\cpu.PCreg1[7] ));
 sg13g2_dfrbp_1 _12847_ (.CLK(net3774),
    .RESET_B(net370),
    .D(_01352_),
    .Q_N(_05762_),
    .Q(\cpu.PCreg1[8] ));
 sg13g2_dfrbp_1 _12848_ (.CLK(net3774),
    .RESET_B(net369),
    .D(_01353_),
    .Q_N(_05761_),
    .Q(\cpu.PCreg1[9] ));
 sg13g2_dfrbp_1 _12849_ (.CLK(net3759),
    .RESET_B(net368),
    .D(_01354_),
    .Q_N(_05760_),
    .Q(\cpu.PCreg1[10] ));
 sg13g2_dfrbp_1 _12850_ (.CLK(net3759),
    .RESET_B(net367),
    .D(_01355_),
    .Q_N(_05759_),
    .Q(\cpu.PCreg1[11] ));
 sg13g2_dfrbp_1 _12851_ (.CLK(net3756),
    .RESET_B(net366),
    .D(_01356_),
    .Q_N(_05758_),
    .Q(\cpu.PCreg1[12] ));
 sg13g2_dfrbp_1 _12852_ (.CLK(net3746),
    .RESET_B(net365),
    .D(_01357_),
    .Q_N(_05757_),
    .Q(\cpu.PCreg1[13] ));
 sg13g2_dfrbp_1 _12853_ (.CLK(net3757),
    .RESET_B(net364),
    .D(_01358_),
    .Q_N(_05756_),
    .Q(\cpu.PCreg1[14] ));
 sg13g2_dfrbp_1 _12854_ (.CLK(net3757),
    .RESET_B(net363),
    .D(_01359_),
    .Q_N(_05755_),
    .Q(\cpu.PCreg1[15] ));
 sg13g2_dfrbp_1 _12855_ (.CLK(net3758),
    .RESET_B(net362),
    .D(_01360_),
    .Q_N(_05754_),
    .Q(\cpu.PCreg1[16] ));
 sg13g2_dfrbp_1 _12856_ (.CLK(net3757),
    .RESET_B(net361),
    .D(_01361_),
    .Q_N(_05753_),
    .Q(\cpu.PCreg1[17] ));
 sg13g2_dfrbp_1 _12857_ (.CLK(net3777),
    .RESET_B(net360),
    .D(_01362_),
    .Q_N(_05752_),
    .Q(\cpu.PCreg1[18] ));
 sg13g2_dfrbp_1 _12858_ (.CLK(net3764),
    .RESET_B(net359),
    .D(_01363_),
    .Q_N(_05751_),
    .Q(\cpu.PCreg1[19] ));
 sg13g2_dfrbp_1 _12859_ (.CLK(net3762),
    .RESET_B(net358),
    .D(_01364_),
    .Q_N(_05750_),
    .Q(\cpu.PCreg1[20] ));
 sg13g2_dfrbp_1 _12860_ (.CLK(net3767),
    .RESET_B(net357),
    .D(_01365_),
    .Q_N(_05749_),
    .Q(\cpu.PCreg1[21] ));
 sg13g2_dfrbp_1 _12861_ (.CLK(net3764),
    .RESET_B(net356),
    .D(_01366_),
    .Q_N(_05748_),
    .Q(\cpu.PCreg1[22] ));
 sg13g2_dfrbp_1 _12862_ (.CLK(net3764),
    .RESET_B(net355),
    .D(_01367_),
    .Q_N(_05747_),
    .Q(\cpu.PCreg1[23] ));
 sg13g2_dfrbp_1 _12863_ (.CLK(net3767),
    .RESET_B(net354),
    .D(_01368_),
    .Q_N(_05746_),
    .Q(\cpu.PCreg1[24] ));
 sg13g2_dfrbp_1 _12864_ (.CLK(net3767),
    .RESET_B(net353),
    .D(_01369_),
    .Q_N(_05745_),
    .Q(\cpu.PCreg1[25] ));
 sg13g2_dfrbp_1 _12865_ (.CLK(net3769),
    .RESET_B(net352),
    .D(_01370_),
    .Q_N(_05744_),
    .Q(\cpu.PCreg1[26] ));
 sg13g2_dfrbp_1 _12866_ (.CLK(net3756),
    .RESET_B(net351),
    .D(_01371_),
    .Q_N(_05743_),
    .Q(\cpu.PCreg1[27] ));
 sg13g2_dfrbp_1 _12867_ (.CLK(net3765),
    .RESET_B(net350),
    .D(_01372_),
    .Q_N(_05742_),
    .Q(\cpu.PCreg1[28] ));
 sg13g2_dfrbp_1 _12868_ (.CLK(net3757),
    .RESET_B(net349),
    .D(_01373_),
    .Q_N(_05741_),
    .Q(\cpu.PCreg1[29] ));
 sg13g2_dfrbp_1 _12869_ (.CLK(net3764),
    .RESET_B(net348),
    .D(_01374_),
    .Q_N(_05740_),
    .Q(\cpu.PCreg1[30] ));
 sg13g2_dfrbp_1 _12870_ (.CLK(net3764),
    .RESET_B(net347),
    .D(_01375_),
    .Q_N(_05739_),
    .Q(\cpu.PCreg1[31] ));
 sg13g2_dfrbp_1 _12871_ (.CLK(net3794),
    .RESET_B(net346),
    .D(_01376_),
    .Q_N(_00123_),
    .Q(\cpu.regs[4][0] ));
 sg13g2_dfrbp_1 _12872_ (.CLK(net3842),
    .RESET_B(net345),
    .D(_01377_),
    .Q_N(_00122_),
    .Q(\cpu.regs[4][1] ));
 sg13g2_dfrbp_1 _12873_ (.CLK(net3792),
    .RESET_B(net344),
    .D(_01378_),
    .Q_N(_00121_),
    .Q(\cpu.regs[4][2] ));
 sg13g2_dfrbp_1 _12874_ (.CLK(net3846),
    .RESET_B(net343),
    .D(_01379_),
    .Q_N(_00120_),
    .Q(\cpu.regs[4][3] ));
 sg13g2_dfrbp_1 _12875_ (.CLK(net3794),
    .RESET_B(net342),
    .D(_01380_),
    .Q_N(_00119_),
    .Q(\cpu.regs[4][4] ));
 sg13g2_dfrbp_1 _12876_ (.CLK(net3863),
    .RESET_B(net341),
    .D(_01381_),
    .Q_N(_00118_),
    .Q(\cpu.regs[4][5] ));
 sg13g2_dfrbp_1 _12877_ (.CLK(net3847),
    .RESET_B(net340),
    .D(_01382_),
    .Q_N(_00117_),
    .Q(\cpu.regs[4][6] ));
 sg13g2_dfrbp_1 _12878_ (.CLK(net3848),
    .RESET_B(net339),
    .D(_01383_),
    .Q_N(_00116_),
    .Q(\cpu.regs[4][7] ));
 sg13g2_dfrbp_1 _12879_ (.CLK(net3845),
    .RESET_B(net338),
    .D(_01384_),
    .Q_N(_00115_),
    .Q(\cpu.regs[4][8] ));
 sg13g2_dfrbp_1 _12880_ (.CLK(net3836),
    .RESET_B(net337),
    .D(_01385_),
    .Q_N(_00114_),
    .Q(\cpu.regs[4][9] ));
 sg13g2_dfrbp_1 _12881_ (.CLK(net3861),
    .RESET_B(net336),
    .D(_01386_),
    .Q_N(_00113_),
    .Q(\cpu.regs[4][10] ));
 sg13g2_dfrbp_1 _12882_ (.CLK(net3856),
    .RESET_B(net335),
    .D(_01387_),
    .Q_N(_00112_),
    .Q(\cpu.regs[4][11] ));
 sg13g2_dfrbp_1 _12883_ (.CLK(net3761),
    .RESET_B(net334),
    .D(_01388_),
    .Q_N(_00111_),
    .Q(\cpu.regs[4][12] ));
 sg13g2_dfrbp_1 _12884_ (.CLK(net3761),
    .RESET_B(net333),
    .D(_01389_),
    .Q_N(_00110_),
    .Q(\cpu.regs[4][13] ));
 sg13g2_dfrbp_1 _12885_ (.CLK(net3834),
    .RESET_B(net332),
    .D(_01390_),
    .Q_N(_00109_),
    .Q(\cpu.regs[4][14] ));
 sg13g2_dfrbp_1 _12886_ (.CLK(net3834),
    .RESET_B(net331),
    .D(_01391_),
    .Q_N(_00108_),
    .Q(\cpu.regs[4][15] ));
 sg13g2_dfrbp_1 _12887_ (.CLK(net3841),
    .RESET_B(net330),
    .D(_01392_),
    .Q_N(_00107_),
    .Q(\cpu.regs[4][16] ));
 sg13g2_dfrbp_1 _12888_ (.CLK(net3853),
    .RESET_B(net329),
    .D(_01393_),
    .Q_N(_00106_),
    .Q(\cpu.regs[4][17] ));
 sg13g2_dfrbp_1 _12889_ (.CLK(net3831),
    .RESET_B(net328),
    .D(_01394_),
    .Q_N(_00105_),
    .Q(\cpu.regs[4][18] ));
 sg13g2_dfrbp_1 _12890_ (.CLK(net3852),
    .RESET_B(net760),
    .D(_01395_),
    .Q_N(_00104_),
    .Q(\cpu.regs[4][19] ));
 sg13g2_dfrbp_1 _12891_ (.CLK(net3761),
    .RESET_B(net759),
    .D(_01396_),
    .Q_N(_00103_),
    .Q(\cpu.regs[4][20] ));
 sg13g2_dfrbp_1 _12892_ (.CLK(net3819),
    .RESET_B(net726),
    .D(_01397_),
    .Q_N(_00102_),
    .Q(\cpu.regs[4][21] ));
 sg13g2_dfrbp_1 _12893_ (.CLK(net3828),
    .RESET_B(net725),
    .D(_01398_),
    .Q_N(_00101_),
    .Q(\cpu.regs[4][22] ));
 sg13g2_dfrbp_1 _12894_ (.CLK(net3821),
    .RESET_B(net724),
    .D(_01399_),
    .Q_N(_00100_),
    .Q(\cpu.regs[4][23] ));
 sg13g2_dfrbp_1 _12895_ (.CLK(net3806),
    .RESET_B(net723),
    .D(_01400_),
    .Q_N(_00099_),
    .Q(\cpu.regs[4][24] ));
 sg13g2_dfrbp_1 _12896_ (.CLK(net3832),
    .RESET_B(net722),
    .D(_01401_),
    .Q_N(_00098_),
    .Q(\cpu.regs[4][25] ));
 sg13g2_dfrbp_1 _12897_ (.CLK(net3800),
    .RESET_B(net721),
    .D(_01402_),
    .Q_N(_00097_),
    .Q(\cpu.regs[4][26] ));
 sg13g2_dfrbp_1 _12898_ (.CLK(net3824),
    .RESET_B(net720),
    .D(_01403_),
    .Q_N(_00096_),
    .Q(\cpu.regs[4][27] ));
 sg13g2_dfrbp_1 _12899_ (.CLK(net3811),
    .RESET_B(net719),
    .D(_01404_),
    .Q_N(_00095_),
    .Q(\cpu.regs[4][28] ));
 sg13g2_dfrbp_1 _12900_ (.CLK(net3827),
    .RESET_B(net718),
    .D(_01405_),
    .Q_N(_00094_),
    .Q(\cpu.regs[4][29] ));
 sg13g2_dfrbp_1 _12901_ (.CLK(net3765),
    .RESET_B(net717),
    .D(_01406_),
    .Q_N(_00093_),
    .Q(\cpu.regs[4][30] ));
 sg13g2_dfrbp_1 _12902_ (.CLK(net3768),
    .RESET_B(net716),
    .D(_01407_),
    .Q_N(_00092_),
    .Q(\cpu.regs[4][31] ));
 sg13g2_dfrbp_1 _12903_ (.CLK(net3792),
    .RESET_B(net715),
    .D(_01408_),
    .Q_N(_00091_),
    .Q(\cpu.regs[3][0] ));
 sg13g2_dfrbp_1 _12904_ (.CLK(net3842),
    .RESET_B(net714),
    .D(_01409_),
    .Q_N(_00090_),
    .Q(\cpu.regs[3][1] ));
 sg13g2_dfrbp_1 _12905_ (.CLK(net3795),
    .RESET_B(net713),
    .D(_01410_),
    .Q_N(_00089_),
    .Q(\cpu.regs[3][2] ));
 sg13g2_dfrbp_1 _12906_ (.CLK(net3846),
    .RESET_B(net712),
    .D(_01411_),
    .Q_N(_00088_),
    .Q(\cpu.regs[3][3] ));
 sg13g2_dfrbp_1 _12907_ (.CLK(net3794),
    .RESET_B(net711),
    .D(_01412_),
    .Q_N(_00087_),
    .Q(\cpu.regs[3][4] ));
 sg13g2_dfrbp_1 _12908_ (.CLK(net3863),
    .RESET_B(net710),
    .D(_01413_),
    .Q_N(_00086_),
    .Q(\cpu.regs[3][5] ));
 sg13g2_dfrbp_1 _12909_ (.CLK(net3843),
    .RESET_B(net709),
    .D(_01414_),
    .Q_N(_00085_),
    .Q(\cpu.regs[3][6] ));
 sg13g2_dfrbp_1 _12910_ (.CLK(net3848),
    .RESET_B(net708),
    .D(_01415_),
    .Q_N(_00084_),
    .Q(\cpu.regs[3][7] ));
 sg13g2_dfrbp_1 _12911_ (.CLK(net3863),
    .RESET_B(net707),
    .D(_01416_),
    .Q_N(_00083_),
    .Q(\cpu.regs[3][8] ));
 sg13g2_dfrbp_1 _12912_ (.CLK(net3836),
    .RESET_B(net706),
    .D(_01417_),
    .Q_N(_00082_),
    .Q(\cpu.regs[3][9] ));
 sg13g2_dfrbp_1 _12913_ (.CLK(net3861),
    .RESET_B(net705),
    .D(_01418_),
    .Q_N(_00081_),
    .Q(\cpu.regs[3][10] ));
 sg13g2_dfrbp_1 _12914_ (.CLK(net3856),
    .RESET_B(net704),
    .D(_01419_),
    .Q_N(_00080_),
    .Q(\cpu.regs[3][11] ));
 sg13g2_dfrbp_1 _12915_ (.CLK(net3799),
    .RESET_B(net703),
    .D(_01420_),
    .Q_N(_00079_),
    .Q(\cpu.regs[3][12] ));
 sg13g2_dfrbp_1 _12916_ (.CLK(net3768),
    .RESET_B(net702),
    .D(_01421_),
    .Q_N(_00078_),
    .Q(\cpu.regs[3][13] ));
 sg13g2_dfrbp_1 _12917_ (.CLK(net3851),
    .RESET_B(net684),
    .D(_01422_),
    .Q_N(_00077_),
    .Q(\cpu.regs[3][14] ));
 sg13g2_dfrbp_1 _12918_ (.CLK(net3811),
    .RESET_B(net538),
    .D(_01423_),
    .Q_N(_00076_),
    .Q(\cpu.regs[3][15] ));
 sg13g2_dfrbp_1 _12919_ (.CLK(net3839),
    .RESET_B(net537),
    .D(_01424_),
    .Q_N(_00075_),
    .Q(\cpu.regs[3][16] ));
 sg13g2_dfrbp_1 _12920_ (.CLK(net3853),
    .RESET_B(net536),
    .D(_01425_),
    .Q_N(_00074_),
    .Q(\cpu.regs[3][17] ));
 sg13g2_dfrbp_1 _12921_ (.CLK(net3831),
    .RESET_B(net534),
    .D(_01426_),
    .Q_N(_00073_),
    .Q(\cpu.regs[3][18] ));
 sg13g2_dfrbp_1 _12922_ (.CLK(net3856),
    .RESET_B(net532),
    .D(_01427_),
    .Q_N(_00072_),
    .Q(\cpu.regs[3][19] ));
 sg13g2_dfrbp_1 _12923_ (.CLK(net3800),
    .RESET_B(net531),
    .D(_01428_),
    .Q_N(_00071_),
    .Q(\cpu.regs[3][20] ));
 sg13g2_dfrbp_1 _12924_ (.CLK(net3818),
    .RESET_B(net529),
    .D(_01429_),
    .Q_N(_00070_),
    .Q(\cpu.regs[3][21] ));
 sg13g2_dfrbp_1 _12925_ (.CLK(net3828),
    .RESET_B(net528),
    .D(_01430_),
    .Q_N(_00069_),
    .Q(\cpu.regs[3][22] ));
 sg13g2_dfrbp_1 _12926_ (.CLK(net3820),
    .RESET_B(net526),
    .D(_01431_),
    .Q_N(_00068_),
    .Q(\cpu.regs[3][23] ));
 sg13g2_dfrbp_1 _12927_ (.CLK(net3810),
    .RESET_B(net525),
    .D(_01432_),
    .Q_N(_00067_),
    .Q(\cpu.regs[3][24] ));
 sg13g2_dfrbp_1 _12928_ (.CLK(net3828),
    .RESET_B(net523),
    .D(_01433_),
    .Q_N(_00066_),
    .Q(\cpu.regs[3][25] ));
 sg13g2_dfrbp_1 _12929_ (.CLK(net3800),
    .RESET_B(net522),
    .D(_01434_),
    .Q_N(_00065_),
    .Q(\cpu.regs[3][26] ));
 sg13g2_dfrbp_1 _12930_ (.CLK(net3825),
    .RESET_B(net520),
    .D(_01435_),
    .Q_N(_00064_),
    .Q(\cpu.regs[3][27] ));
 sg13g2_dfrbp_1 _12931_ (.CLK(net3811),
    .RESET_B(net519),
    .D(_01436_),
    .Q_N(_00063_),
    .Q(\cpu.regs[3][28] ));
 sg13g2_dfrbp_1 _12932_ (.CLK(net3811),
    .RESET_B(net517),
    .D(_01437_),
    .Q_N(_00062_),
    .Q(\cpu.regs[3][29] ));
 sg13g2_dfrbp_1 _12933_ (.CLK(net3767),
    .RESET_B(net516),
    .D(_01438_),
    .Q_N(_00061_),
    .Q(\cpu.regs[3][30] ));
 sg13g2_dfrbp_1 _12934_ (.CLK(net3799),
    .RESET_B(net514),
    .D(_01439_),
    .Q_N(_00060_),
    .Q(\cpu.regs[3][31] ));
 sg13g2_dfrbp_1 _12935_ (.CLK(net3920),
    .RESET_B(net3714),
    .D(_00691_),
    .Q_N(\uart0.urxsh[0] ),
    .Q(_00581_));
 sg13g2_dfrbp_1 _12936_ (.CLK(clknet_2_0__leaf_jclk_regs),
    .RESET_B(net511),
    .D(_01440_),
    .Q_N(_05738_),
    .Q(\xdi[16] ));
 sg13g2_dfrbp_1 _12937_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net510),
    .D(net911),
    .Q_N(_05737_),
    .Q(\xdi[17] ));
 sg13g2_dfrbp_1 _12938_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net508),
    .D(net924),
    .Q_N(_05736_),
    .Q(\xdi[18] ));
 sg13g2_dfrbp_1 _12939_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net507),
    .D(_01443_),
    .Q_N(_05735_),
    .Q(\xdi[19] ));
 sg13g2_dfrbp_1 _12940_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net505),
    .D(_01444_),
    .Q_N(_05734_),
    .Q(\xdi[20] ));
 sg13g2_dfrbp_1 _12941_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net504),
    .D(net894),
    .Q_N(_05733_),
    .Q(\xdi[21] ));
 sg13g2_dfrbp_1 _12942_ (.CLK(clknet_2_3__leaf_jclk_regs),
    .RESET_B(net502),
    .D(_01446_),
    .Q_N(_05732_),
    .Q(\xdi[22] ));
 sg13g2_dfrbp_1 _12943_ (.CLK(clknet_2_1__leaf_jclk_regs),
    .RESET_B(net728),
    .D(net913),
    .Q_N(_06039_),
    .Q(\xdi[23] ));
 sg13g2_dfrbp_1 _12944_ (.CLK(net3785),
    .RESET_B(net3721),
    .D(_00013_),
    .Q_N(_00546_),
    .Q(\cpu.opvalid ));
 sg13g2_dfrbp_1 _12945_ (.CLK(net3781),
    .RESET_B(net729),
    .D(\cdi[0] ),
    .Q_N(_06040_),
    .Q(\cpu.IR[0] ));
 sg13g2_dfrbp_1 _12946_ (.CLK(net3781),
    .RESET_B(net730),
    .D(\cdi[1] ),
    .Q_N(_06041_),
    .Q(\cpu.IR[1] ));
 sg13g2_dfrbp_1 _12947_ (.CLK(net3781),
    .RESET_B(net731),
    .D(\cdi[2] ),
    .Q_N(_06042_),
    .Q(\cpu.IR[2] ));
 sg13g2_dfrbp_1 _12948_ (.CLK(net3781),
    .RESET_B(net732),
    .D(\cdi[3] ),
    .Q_N(_06043_),
    .Q(\cpu.IR[3] ));
 sg13g2_dfrbp_1 _12949_ (.CLK(net3782),
    .RESET_B(net733),
    .D(\cdi[4] ),
    .Q_N(_06044_),
    .Q(\cpu.IR[4] ));
 sg13g2_dfrbp_1 _12950_ (.CLK(net3782),
    .RESET_B(net734),
    .D(\cdi[5] ),
    .Q_N(_06045_),
    .Q(\cpu.IR[5] ));
 sg13g2_dfrbp_1 _12951_ (.CLK(net3783),
    .RESET_B(net735),
    .D(\cdi[6] ),
    .Q_N(_00547_),
    .Q(\cpu.IR[6] ));
 sg13g2_dfrbp_1 _12952_ (.CLK(net3781),
    .RESET_B(net736),
    .D(\cdi[7] ),
    .Q_N(_06046_),
    .Q(\cpu.Bimm[11] ));
 sg13g2_dfrbp_1 _12953_ (.CLK(net3783),
    .RESET_B(net737),
    .D(\cdi[8] ),
    .Q_N(_00548_),
    .Q(\cpu.Bimm[1] ));
 sg13g2_dfrbp_1 _12954_ (.CLK(net3839),
    .RESET_B(net738),
    .D(\cdi[9] ),
    .Q_N(_00549_),
    .Q(\cpu.Bimm[2] ));
 sg13g2_dfrbp_1 _12955_ (.CLK(net3839),
    .RESET_B(net739),
    .D(\cdi[10] ),
    .Q_N(_00550_),
    .Q(\cpu.Bimm[3] ));
 sg13g2_dfrbp_1 _12956_ (.CLK(net3784),
    .RESET_B(net740),
    .D(\cdi[11] ),
    .Q_N(_00551_),
    .Q(\cpu.Bimm[4] ));
 sg13g2_dfrbp_1 _12957_ (.CLK(net3782),
    .RESET_B(net741),
    .D(\cdi[12] ),
    .Q_N(_06047_),
    .Q(\cpu.IR[12] ));
 sg13g2_dfrbp_1 _12958_ (.CLK(net3759),
    .RESET_B(net742),
    .D(\cdi[13] ),
    .Q_N(_06048_),
    .Q(\cpu.IR[13] ));
 sg13g2_dfrbp_1 _12959_ (.CLK(net3785),
    .RESET_B(net743),
    .D(\cdi[14] ),
    .Q_N(_00552_),
    .Q(\cpu.IR[14] ));
 sg13g2_dfrbp_1 _12960_ (.CLK(net3782),
    .RESET_B(net744),
    .D(\cdi[15] ),
    .Q_N(_06049_),
    .Q(\cpu.IR[15] ));
 sg13g2_dfrbp_1 _12961_ (.CLK(net3783),
    .RESET_B(net745),
    .D(\cdi[16] ),
    .Q_N(_06050_),
    .Q(\cpu.IR[16] ));
 sg13g2_dfrbp_1 _12962_ (.CLK(net3839),
    .RESET_B(net746),
    .D(\cdi[17] ),
    .Q_N(_06051_),
    .Q(\cpu.IR[17] ));
 sg13g2_dfrbp_1 _12963_ (.CLK(net3809),
    .RESET_B(net747),
    .D(\cdi[18] ),
    .Q_N(_06052_),
    .Q(\cpu.IR[18] ));
 sg13g2_dfrbp_1 _12964_ (.CLK(net3777),
    .RESET_B(net748),
    .D(\cdi[19] ),
    .Q_N(_06053_),
    .Q(\cpu.IR[19] ));
 sg13g2_dfrbp_1 _12965_ (.CLK(net3774),
    .RESET_B(net749),
    .D(\cdi[20] ),
    .Q_N(_06054_),
    .Q(\cpu.IR[20] ));
 sg13g2_dfrbp_1 _12966_ (.CLK(net3783),
    .RESET_B(net750),
    .D(\cdi[21] ),
    .Q_N(_00553_),
    .Q(\cpu.IR[21] ));
 sg13g2_dfrbp_1 _12967_ (.CLK(net3784),
    .RESET_B(net751),
    .D(\cdi[22] ),
    .Q_N(_00554_),
    .Q(\cpu.IR[22] ));
 sg13g2_dfrbp_1 _12968_ (.CLK(net3784),
    .RESET_B(net752),
    .D(\cdi[23] ),
    .Q_N(_00555_),
    .Q(\cpu.IR[23] ));
 sg13g2_dfrbp_1 _12969_ (.CLK(net3784),
    .RESET_B(net753),
    .D(\cdi[24] ),
    .Q_N(_00556_),
    .Q(\cpu.IR[24] ));
 sg13g2_dfrbp_1 _12970_ (.CLK(net3784),
    .RESET_B(net754),
    .D(\cdi[25] ),
    .Q_N(_00557_),
    .Q(\cpu.Bimm[5] ));
 sg13g2_dfrbp_1 _12971_ (.CLK(net3785),
    .RESET_B(net755),
    .D(\cdi[26] ),
    .Q_N(_00558_),
    .Q(\cpu.Bimm[6] ));
 sg13g2_dfrbp_1 _12972_ (.CLK(net3785),
    .RESET_B(net756),
    .D(\cdi[27] ),
    .Q_N(_00559_),
    .Q(\cpu.Bimm[7] ));
 sg13g2_dfrbp_1 _12973_ (.CLK(net3782),
    .RESET_B(net757),
    .D(\cdi[28] ),
    .Q_N(_00560_),
    .Q(\cpu.Bimm[8] ));
 sg13g2_dfrbp_1 _12974_ (.CLK(net3774),
    .RESET_B(net758),
    .D(\cdi[29] ),
    .Q_N(_00561_),
    .Q(\cpu.Bimm[9] ));
 sg13g2_dfrbp_1 _12975_ (.CLK(net3774),
    .RESET_B(net788),
    .D(\cdi[30] ),
    .Q_N(_00562_),
    .Q(\cpu.Bimm[10] ));
 sg13g2_dfrbp_1 _12976_ (.CLK(net3775),
    .RESET_B(net501),
    .D(\cdi[31] ),
    .Q_N(_00059_),
    .Q(\cpu.Bimm[12] ));
 sg13g2_dfrbp_1 _12977_ (.CLK(net3792),
    .RESET_B(net3721),
    .D(_01448_),
    .Q_N(_05731_),
    .Q(\cpu.PCreg0[2] ));
 sg13g2_dfrbp_1 _12978_ (.CLK(net3783),
    .RESET_B(net3721),
    .D(_01449_),
    .Q_N(_05730_),
    .Q(\cpu.PCreg0[3] ));
 sg13g2_dfrbp_1 _12979_ (.CLK(net3781),
    .RESET_B(net3721),
    .D(_01450_),
    .Q_N(_05729_),
    .Q(\cpu.PCreg0[4] ));
 sg13g2_dfrbp_1 _12980_ (.CLK(net3781),
    .RESET_B(net3721),
    .D(_01451_),
    .Q_N(_05728_),
    .Q(\cpu.PCreg0[5] ));
 sg13g2_dfrbp_1 _12981_ (.CLK(net3783),
    .RESET_B(net3721),
    .D(_01452_),
    .Q_N(_05727_),
    .Q(\cpu.PCreg0[6] ));
 sg13g2_dfrbp_1 _12982_ (.CLK(net3774),
    .RESET_B(net3712),
    .D(_01453_),
    .Q_N(_05726_),
    .Q(\cpu.PCreg0[7] ));
 sg13g2_dfrbp_1 _12983_ (.CLK(net3782),
    .RESET_B(net3711),
    .D(_01454_),
    .Q_N(_05725_),
    .Q(\cpu.PCreg0[8] ));
 sg13g2_dfrbp_1 _12984_ (.CLK(net3775),
    .RESET_B(net3712),
    .D(_01455_),
    .Q_N(_05724_),
    .Q(\cpu.PCreg0[9] ));
 sg13g2_dfrbp_1 _12985_ (.CLK(net3774),
    .RESET_B(net3711),
    .D(_01456_),
    .Q_N(_05723_),
    .Q(\cpu.PCreg0[10] ));
 sg13g2_dfrbp_1 _12986_ (.CLK(net3774),
    .RESET_B(net3711),
    .D(_01457_),
    .Q_N(_05722_),
    .Q(\cpu.PCreg0[11] ));
 sg13g2_dfrbp_1 _12987_ (.CLK(net3772),
    .RESET_B(net3711),
    .D(_01458_),
    .Q_N(_05721_),
    .Q(\cpu.PCreg0[12] ));
 sg13g2_dfrbp_1 _12988_ (.CLK(net3772),
    .RESET_B(net3708),
    .D(_01459_),
    .Q_N(_05720_),
    .Q(\cpu.PCreg0[13] ));
 sg13g2_dfrbp_1 _12989_ (.CLK(net3772),
    .RESET_B(net3711),
    .D(_01460_),
    .Q_N(_05719_),
    .Q(\cpu.PCreg0[14] ));
 sg13g2_dfrbp_1 _12990_ (.CLK(net3772),
    .RESET_B(net3711),
    .D(_01461_),
    .Q_N(_05718_),
    .Q(\cpu.PCreg0[15] ));
 sg13g2_dfrbp_1 _12991_ (.CLK(net3773),
    .RESET_B(net3708),
    .D(_01462_),
    .Q_N(_05717_),
    .Q(\cpu.PCreg0[16] ));
 sg13g2_dfrbp_1 _12992_ (.CLK(net3772),
    .RESET_B(net3708),
    .D(_01463_),
    .Q_N(_05716_),
    .Q(\cpu.PCreg0[17] ));
 sg13g2_dfrbp_1 _12993_ (.CLK(net3777),
    .RESET_B(net3710),
    .D(_01464_),
    .Q_N(_05715_),
    .Q(\cpu.PCreg0[18] ));
 sg13g2_dfrbp_1 _12994_ (.CLK(net3770),
    .RESET_B(net3709),
    .D(_01465_),
    .Q_N(_05714_),
    .Q(\cpu.PCreg0[19] ));
 sg13g2_dfrbp_1 _12995_ (.CLK(net3765),
    .RESET_B(net3707),
    .D(_01466_),
    .Q_N(_05713_),
    .Q(\cpu.PCreg0[20] ));
 sg13g2_dfrbp_1 _12996_ (.CLK(net3768),
    .RESET_B(net3709),
    .D(_01467_),
    .Q_N(_05712_),
    .Q(\cpu.PCreg0[21] ));
 sg13g2_dfrbp_1 _12997_ (.CLK(net3770),
    .RESET_B(net3709),
    .D(_01468_),
    .Q_N(_05711_),
    .Q(\cpu.PCreg0[22] ));
 sg13g2_dfrbp_1 _12998_ (.CLK(net3770),
    .RESET_B(net3709),
    .D(_01469_),
    .Q_N(_05710_),
    .Q(\cpu.PCreg0[23] ));
 sg13g2_dfrbp_1 _12999_ (.CLK(net3770),
    .RESET_B(net3709),
    .D(_01470_),
    .Q_N(_05709_),
    .Q(\cpu.PCreg0[24] ));
 sg13g2_dfrbp_1 _13000_ (.CLK(net3769),
    .RESET_B(net3709),
    .D(_01471_),
    .Q_N(_05708_),
    .Q(\cpu.PCreg0[25] ));
 sg13g2_dfrbp_1 _13001_ (.CLK(net3770),
    .RESET_B(net3709),
    .D(_01472_),
    .Q_N(_05707_),
    .Q(\cpu.PCreg0[26] ));
 sg13g2_dfrbp_1 _13002_ (.CLK(net3772),
    .RESET_B(net3710),
    .D(_01473_),
    .Q_N(_05706_),
    .Q(\cpu.PCreg0[27] ));
 sg13g2_dfrbp_1 _13003_ (.CLK(net3765),
    .RESET_B(net3709),
    .D(_01474_),
    .Q_N(_05705_),
    .Q(\cpu.PCreg0[28] ));
 sg13g2_dfrbp_1 _13004_ (.CLK(net3773),
    .RESET_B(net3708),
    .D(_01475_),
    .Q_N(_05704_),
    .Q(\cpu.PCreg0[29] ));
 sg13g2_dfrbp_1 _13005_ (.CLK(net3764),
    .RESET_B(net3708),
    .D(_01476_),
    .Q_N(_05703_),
    .Q(\cpu.PCreg0[30] ));
 sg13g2_dfrbp_1 _13006_ (.CLK(net3764),
    .RESET_B(net3707),
    .D(_01477_),
    .Q_N(_06055_),
    .Q(\cpu.PCreg0[31] ));
 sg13g2_dfrbp_1 _13007_ (.CLK(net3796),
    .RESET_B(net789),
    .D(\cpu.PC[2] ),
    .Q_N(_00563_),
    .Q(\cpu.PCci[2] ));
 sg13g2_dfrbp_1 _13008_ (.CLK(net3784),
    .RESET_B(net790),
    .D(\cpu.PC[3] ),
    .Q_N(_00564_),
    .Q(\cpu.PCci[3] ));
 sg13g2_dfrbp_1 _13009_ (.CLK(net3783),
    .RESET_B(net791),
    .D(\cpu.PC[4] ),
    .Q_N(_00565_),
    .Q(\cpu.PCci[4] ));
 sg13g2_dfrbp_1 _13010_ (.CLK(net3783),
    .RESET_B(net792),
    .D(\cpu.PC[5] ),
    .Q_N(_06056_),
    .Q(\cpu.PCci[5] ));
 sg13g2_dfrbp_1 _13011_ (.CLK(net3785),
    .RESET_B(net793),
    .D(\cpu.PC[6] ),
    .Q_N(_00566_),
    .Q(\cpu.PCci[6] ));
 sg13g2_dfrbp_1 _13012_ (.CLK(net3785),
    .RESET_B(net794),
    .D(\cpu.PC[7] ),
    .Q_N(_06057_),
    .Q(\cpu.PCci[7] ));
 sg13g2_dfrbp_1 _13013_ (.CLK(net3777),
    .RESET_B(net795),
    .D(\cpu.PC[8] ),
    .Q_N(_00567_),
    .Q(\cpu.PCci[8] ));
 sg13g2_dfrbp_1 _13014_ (.CLK(net3778),
    .RESET_B(net796),
    .D(\cpu.PC[9] ),
    .Q_N(_06058_),
    .Q(\cpu.PCci[9] ));
 sg13g2_dfrbp_1 _13015_ (.CLK(net3777),
    .RESET_B(net797),
    .D(\cpu.PC[10] ),
    .Q_N(_00568_),
    .Q(\cpu.PCci[10] ));
 sg13g2_dfrbp_1 _13016_ (.CLK(net3777),
    .RESET_B(net798),
    .D(\cpu.PC[11] ),
    .Q_N(_06059_),
    .Q(\cpu.PCci[11] ));
 sg13g2_dfrbp_1 _13017_ (.CLK(net3777),
    .RESET_B(net799),
    .D(\cpu.PC[12] ),
    .Q_N(_00569_),
    .Q(\cpu.PCci[12] ));
 sg13g2_dfrbp_1 _13018_ (.CLK(net3775),
    .RESET_B(net800),
    .D(\cpu.PC[13] ),
    .Q_N(_06060_),
    .Q(\cpu.PCci[13] ));
 sg13g2_dfrbp_1 _13019_ (.CLK(net3775),
    .RESET_B(net801),
    .D(\cpu.PC[14] ),
    .Q_N(_06061_),
    .Q(\cpu.PCci[14] ));
 sg13g2_dfrbp_1 _13020_ (.CLK(net3773),
    .RESET_B(net802),
    .D(\cpu.PC[15] ),
    .Q_N(_06062_),
    .Q(\cpu.PCci[15] ));
 sg13g2_dfrbp_1 _13021_ (.CLK(net3772),
    .RESET_B(net803),
    .D(\cpu.PC[16] ),
    .Q_N(_06063_),
    .Q(\cpu.PCci[16] ));
 sg13g2_dfrbp_1 _13022_ (.CLK(net3777),
    .RESET_B(net804),
    .D(\cpu.PC[17] ),
    .Q_N(_06064_),
    .Q(\cpu.PCci[17] ));
 sg13g2_dfrbp_1 _13023_ (.CLK(net3771),
    .RESET_B(net805),
    .D(\cpu.PC[18] ),
    .Q_N(_06065_),
    .Q(\cpu.PCci[18] ));
 sg13g2_dfrbp_1 _13024_ (.CLK(net3770),
    .RESET_B(net806),
    .D(\cpu.PC[19] ),
    .Q_N(_00570_),
    .Q(\cpu.PCci[19] ));
 sg13g2_dfrbp_1 _13025_ (.CLK(net3802),
    .RESET_B(net807),
    .D(\cpu.PC[20] ),
    .Q_N(_06066_),
    .Q(\cpu.PCci[20] ));
 sg13g2_dfrbp_1 _13026_ (.CLK(net3799),
    .RESET_B(net808),
    .D(\cpu.PC[21] ),
    .Q_N(_06067_),
    .Q(\cpu.PCci[21] ));
 sg13g2_dfrbp_1 _13027_ (.CLK(net3801),
    .RESET_B(net809),
    .D(\cpu.PC[22] ),
    .Q_N(_06068_),
    .Q(\cpu.PCci[22] ));
 sg13g2_dfrbp_1 _13028_ (.CLK(net3799),
    .RESET_B(net810),
    .D(\cpu.PC[23] ),
    .Q_N(_00571_),
    .Q(\cpu.PCci[23] ));
 sg13g2_dfrbp_1 _13029_ (.CLK(net3768),
    .RESET_B(net811),
    .D(\cpu.PC[24] ),
    .Q_N(_06069_),
    .Q(\cpu.PCci[24] ));
 sg13g2_dfrbp_1 _13030_ (.CLK(net3768),
    .RESET_B(net812),
    .D(\cpu.PC[25] ),
    .Q_N(_06070_),
    .Q(\cpu.PCci[25] ));
 sg13g2_dfrbp_1 _13031_ (.CLK(net3771),
    .RESET_B(net813),
    .D(\cpu.PC[26] ),
    .Q_N(_06071_),
    .Q(\cpu.PCci[26] ));
 sg13g2_dfrbp_1 _13032_ (.CLK(net3770),
    .RESET_B(net814),
    .D(\cpu.PC[27] ),
    .Q_N(_06072_),
    .Q(\cpu.PCci[27] ));
 sg13g2_dfrbp_1 _13033_ (.CLK(net3770),
    .RESET_B(net815),
    .D(\cpu.PC[28] ),
    .Q_N(_06073_),
    .Q(\cpu.PCci[28] ));
 sg13g2_dfrbp_1 _13034_ (.CLK(net3772),
    .RESET_B(net816),
    .D(\cpu.PC[29] ),
    .Q_N(_06074_),
    .Q(\cpu.PCci[29] ));
 sg13g2_dfrbp_1 _13035_ (.CLK(net3773),
    .RESET_B(net817),
    .D(\cpu.PC[30] ),
    .Q_N(_06075_),
    .Q(\cpu.PCci[30] ));
 sg13g2_dfrbp_1 _13036_ (.CLK(net3764),
    .RESET_B(net818),
    .D(\cpu.PC[31] ),
    .Q_N(_06076_),
    .Q(\cpu.PCci[31] ));
 sg13g2_dfrbp_1 _13037_ (.CLK(net3782),
    .RESET_B(net3711),
    .D(_00012_),
    .Q_N(_06077_),
    .Q(\cpu.mmode ));
 sg13g2_dfrbp_1 _13038_ (.CLK(net3782),
    .RESET_B(net3711),
    .D(_00014_),
    .Q_N(_05702_),
    .Q(\cpu.q0 ));
 sg13g2_dfrbp_1 _13039_ (.CLK(net3750),
    .RESET_B(net484),
    .D(_01478_),
    .Q_N(_05701_),
    .Q(\irqvect[3][0] ));
 sg13g2_dfrbp_1 _13040_ (.CLK(net3753),
    .RESET_B(net483),
    .D(_01479_),
    .Q_N(_05700_),
    .Q(\irqvect[3][1] ));
 sg13g2_dfrbp_1 _13041_ (.CLK(net3751),
    .RESET_B(net480),
    .D(_01480_),
    .Q_N(_05699_),
    .Q(\irqvect[3][2] ));
 sg13g2_dfrbp_1 _13042_ (.CLK(net3753),
    .RESET_B(net479),
    .D(_01481_),
    .Q_N(_05698_),
    .Q(\irqvect[3][3] ));
 sg13g2_dfrbp_1 _13043_ (.CLK(net3779),
    .RESET_B(net477),
    .D(_01482_),
    .Q_N(_05697_),
    .Q(\irqvect[3][4] ));
 sg13g2_dfrbp_1 _13044_ (.CLK(net3754),
    .RESET_B(net476),
    .D(_01483_),
    .Q_N(_05696_),
    .Q(\irqvect[3][5] ));
 sg13g2_dfrbp_1 _13045_ (.CLK(net3754),
    .RESET_B(net474),
    .D(_01484_),
    .Q_N(_05695_),
    .Q(\irqvect[3][6] ));
 sg13g2_dfrbp_1 _13046_ (.CLK(net3754),
    .RESET_B(net473),
    .D(_01485_),
    .Q_N(_05694_),
    .Q(\irqvect[3][7] ));
 sg13g2_dfrbp_1 _13047_ (.CLK(net3759),
    .RESET_B(net471),
    .D(_01486_),
    .Q_N(_05693_),
    .Q(\irqvect[3][8] ));
 sg13g2_dfrbp_1 _13048_ (.CLK(net3747),
    .RESET_B(net470),
    .D(_01487_),
    .Q_N(_05692_),
    .Q(\irqvect[3][9] ));
 sg13g2_dfrbp_1 _13049_ (.CLK(net3752),
    .RESET_B(net468),
    .D(_01488_),
    .Q_N(_05691_),
    .Q(\irqvect[3][10] ));
 sg13g2_dfrbp_1 _13050_ (.CLK(net3742),
    .RESET_B(net466),
    .D(_01489_),
    .Q_N(_05690_),
    .Q(\irqvect[3][11] ));
 sg13g2_dfrbp_1 _13051_ (.CLK(net3745),
    .RESET_B(net464),
    .D(_01490_),
    .Q_N(_05689_),
    .Q(\irqvect[3][12] ));
 sg13g2_dfrbp_1 _13052_ (.CLK(net3757),
    .RESET_B(net462),
    .D(_01491_),
    .Q_N(_05688_),
    .Q(\irqvect[3][13] ));
 sg13g2_dfrbp_1 _13053_ (.CLK(net3752),
    .RESET_B(net460),
    .D(_01492_),
    .Q_N(_05687_),
    .Q(\irqvect[3][14] ));
 sg13g2_dfrbp_1 _13054_ (.CLK(net3751),
    .RESET_B(net458),
    .D(_01493_),
    .Q_N(_05686_),
    .Q(\irqvect[3][15] ));
 sg13g2_dfrbp_1 _13055_ (.CLK(net3750),
    .RESET_B(net456),
    .D(_01494_),
    .Q_N(_05685_),
    .Q(\irqvect[3][16] ));
 sg13g2_dfrbp_1 _13056_ (.CLK(net3746),
    .RESET_B(net454),
    .D(_01495_),
    .Q_N(_05684_),
    .Q(\irqvect[3][17] ));
 sg13g2_dfrbp_1 _13057_ (.CLK(net3744),
    .RESET_B(net452),
    .D(_01496_),
    .Q_N(_05683_),
    .Q(\irqvect[3][18] ));
 sg13g2_dfrbp_1 _13058_ (.CLK(net3749),
    .RESET_B(net450),
    .D(_01497_),
    .Q_N(_05682_),
    .Q(\irqvect[3][19] ));
 sg13g2_dfrbp_1 _13059_ (.CLK(net3745),
    .RESET_B(net448),
    .D(_01498_),
    .Q_N(_05681_),
    .Q(\irqvect[3][20] ));
 sg13g2_dfrbp_1 _13060_ (.CLK(net3747),
    .RESET_B(net446),
    .D(_01499_),
    .Q_N(_05680_),
    .Q(\irqvect[3][21] ));
 sg13g2_dfrbp_1 _13061_ (.CLK(net3743),
    .RESET_B(net444),
    .D(_01500_),
    .Q_N(_05679_),
    .Q(\irqvect[3][22] ));
 sg13g2_dfrbp_1 _13062_ (.CLK(net3762),
    .RESET_B(net442),
    .D(_01501_),
    .Q_N(_05678_),
    .Q(\irqvect[3][23] ));
 sg13g2_dfrbp_1 _13063_ (.CLK(net3762),
    .RESET_B(net440),
    .D(_01502_),
    .Q_N(_05677_),
    .Q(\irqvect[3][24] ));
 sg13g2_dfrbp_1 _13064_ (.CLK(net3757),
    .RESET_B(net438),
    .D(_01503_),
    .Q_N(_05676_),
    .Q(\irqvect[3][25] ));
 sg13g2_dfrbp_1 _13065_ (.CLK(net3744),
    .RESET_B(net436),
    .D(_01504_),
    .Q_N(_05675_),
    .Q(\irqvect[3][26] ));
 sg13g2_dfrbp_1 _13066_ (.CLK(net3756),
    .RESET_B(net434),
    .D(_01505_),
    .Q_N(_05674_),
    .Q(\irqvect[3][27] ));
 sg13g2_dfrbp_1 _13067_ (.CLK(net3741),
    .RESET_B(net432),
    .D(_01506_),
    .Q_N(_05673_),
    .Q(\irqvect[3][28] ));
 sg13g2_dfrbp_1 _13068_ (.CLK(net3740),
    .RESET_B(net430),
    .D(_01507_),
    .Q_N(_05672_),
    .Q(\irqvect[3][29] ));
 sg13g2_dfrbp_1 _13069_ (.CLK(net3913),
    .RESET_B(net3714),
    .D(_01508_),
    .Q_N(\uart0.urxsh[1] ),
    .Q(_00582_));
 sg13g2_dfrbp_1 _13070_ (.CLK(net3913),
    .RESET_B(net3714),
    .D(_01509_),
    .Q_N(\uart0.urxsh[2] ),
    .Q(_00583_));
 sg13g2_dfrbp_1 _13071_ (.CLK(net3912),
    .RESET_B(net3713),
    .D(_01510_),
    .Q_N(\uart0.urxsh[3] ),
    .Q(_00584_));
 sg13g2_dfrbp_1 _13072_ (.CLK(net3912),
    .RESET_B(net3713),
    .D(_01511_),
    .Q_N(\uart0.urxsh[4] ),
    .Q(_00585_));
 sg13g2_dfrbp_1 _13073_ (.CLK(net3911),
    .RESET_B(net3714),
    .D(_01512_),
    .Q_N(\uart0.urxsh[5] ),
    .Q(_00586_));
 sg13g2_dfrbp_1 _13074_ (.CLK(net3911),
    .RESET_B(net3713),
    .D(_01513_),
    .Q_N(\uart0.urxsh[6] ),
    .Q(_00587_));
 sg13g2_dfrbp_1 _13075_ (.CLK(net3911),
    .RESET_B(net3714),
    .D(_01514_),
    .Q_N(\uart0.urxsh[7] ),
    .Q(_00588_));
 sg13g2_dfrbp_1 _13076_ (.CLK(net3911),
    .RESET_B(net3713),
    .D(_01515_),
    .Q_N(\uart0.urxsh[8] ),
    .Q(_00589_));
 sg13g2_dfrbp_1 _13077_ (.CLK(net3911),
    .RESET_B(net3713),
    .D(_01516_),
    .Q_N(\uart0.urxsh[9] ),
    .Q(_00590_));
 sg13g2_dfrbp_1 _13078_ (.CLK(net3913),
    .RESET_B(net3706),
    .D(_00015_),
    .Q_N(_05671_),
    .Q(\uart0.rxdiv[0] ));
 sg13g2_dfrbp_1 _13079_ (.CLK(net3913),
    .RESET_B(net3706),
    .D(_00016_),
    .Q_N(_05670_),
    .Q(\uart0.rxdiv[1] ));
 sg13g2_dfrbp_1 _13080_ (.CLK(net3913),
    .RESET_B(net3713),
    .D(_00017_),
    .Q_N(_05669_),
    .Q(\uart0.rxdiv[2] ));
 sg13g2_dfrbp_1 _13081_ (.CLK(net3911),
    .RESET_B(net3713),
    .D(_00018_),
    .Q_N(_05668_),
    .Q(\uart0.rxdiv[3] ));
 sg13g2_dfrbp_1 _13082_ (.CLK(net3911),
    .RESET_B(net3713),
    .D(_00019_),
    .Q_N(_05667_),
    .Q(\uart0.rxdiv[4] ));
 sg13g2_dfrbp_1 _13083_ (.CLK(net3913),
    .RESET_B(net3706),
    .D(_00020_),
    .Q_N(_05666_),
    .Q(\uart0.rxdiv[5] ));
 sg13g2_dfrbp_1 _13084_ (.CLK(net3916),
    .RESET_B(net3716),
    .D(_01517_),
    .Q_N(_05665_),
    .Q(\uart0.txbitcnt[0] ));
 sg13g2_dfrbp_1 _13085_ (.CLK(net3915),
    .RESET_B(net3716),
    .D(_01518_),
    .Q_N(_05664_),
    .Q(\uart0.txbitcnt[1] ));
 sg13g2_dfrbp_1 _13086_ (.CLK(net3915),
    .RESET_B(net3716),
    .D(_01519_),
    .Q_N(_05663_),
    .Q(\uart0.txbitcnt[2] ));
 sg13g2_dfrbp_1 _13087_ (.CLK(net3915),
    .RESET_B(net3716),
    .D(_01520_),
    .Q_N(_05662_),
    .Q(\uart0.txbitcnt[3] ));
 sg13g2_dfrbp_1 _13088_ (.CLK(net3914),
    .RESET_B(net416),
    .D(_01521_),
    .Q_N(_05661_),
    .Q(\uart0.q[0] ));
 sg13g2_dfrbp_1 _13089_ (.CLK(net3914),
    .RESET_B(net412),
    .D(_01522_),
    .Q_N(_05660_),
    .Q(\uart0.q[1] ));
 sg13g2_dfrbp_1 _13090_ (.CLK(net3914),
    .RESET_B(net407),
    .D(_01523_),
    .Q_N(_05659_),
    .Q(\uart0.q[2] ));
 sg13g2_dfrbp_1 _13091_ (.CLK(net3911),
    .RESET_B(net404),
    .D(_01524_),
    .Q_N(_05658_),
    .Q(\uart0.q[3] ));
 sg13g2_dfrbp_1 _13092_ (.CLK(net3912),
    .RESET_B(net399),
    .D(_01525_),
    .Q_N(_05657_),
    .Q(\uart0.q[4] ));
 sg13g2_dfrbp_1 _13093_ (.CLK(net3912),
    .RESET_B(net395),
    .D(_01526_),
    .Q_N(_05656_),
    .Q(\uart0.q[5] ));
 sg13g2_dfrbp_1 _13094_ (.CLK(net3915),
    .RESET_B(net391),
    .D(_01527_),
    .Q_N(_05655_),
    .Q(\uart0.q[6] ));
 sg13g2_dfrbp_1 _13095_ (.CLK(net3915),
    .RESET_B(net387),
    .D(_01528_),
    .Q_N(_05654_),
    .Q(\uart0.q[7] ));
 sg13g2_dfrbp_1 _13096_ (.CLK(net3915),
    .RESET_B(net383),
    .D(_01529_),
    .Q_N(_05653_),
    .Q(\uart0.urxbuffer[8] ));
 sg13g2_dfrbp_1 _13097_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(rxd),
    .Q_N(_05652_),
    .Q(\uart0.rxreg[0] ));
 sg13g2_dfrbp_1 _13098_ (.CLK(net3915),
    .RESET_B(net3716),
    .D(\uart0.rxreg[0] ),
    .Q_N(_05651_),
    .Q(\uart0.rxreg[1] ));
 sg13g2_dfrbp_1 _13099_ (.CLK(net3914),
    .RESET_B(net3719),
    .D(_01530_),
    .Q_N(_05650_),
    .Q(\uart0.rxvalid ));
 sg13g2_dfrbp_1 _13100_ (.CLK(net3914),
    .RESET_B(net3714),
    .D(_01531_),
    .Q_N(_05649_),
    .Q(\uart0.rxoverr ));
 sg13g2_dfrbp_1 _13101_ (.CLK(_00692_),
    .RESET_B(net410),
    .D(_01532_),
    .Q_N(_05648_),
    .Q(\jtag0.irsh[0] ));
 sg13g2_dfrbp_1 _13102_ (.CLK(_00693_),
    .RESET_B(net401),
    .D(_01533_),
    .Q_N(_05647_),
    .Q(\jtag0.irsh[1] ));
 sg13g2_dfrbp_1 _13103_ (.CLK(_00694_),
    .RESET_B(net393),
    .D(_01534_),
    .Q_N(_05646_),
    .Q(\jtag0.irsh[2] ));
 sg13g2_dfrbp_1 _13104_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00021_),
    .Q_N(_05645_),
    .Q(\uart0.txdiv[0] ));
 sg13g2_dfrbp_1 _13105_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00022_),
    .Q_N(_05644_),
    .Q(\uart0.txdiv[1] ));
 sg13g2_dfrbp_1 _13106_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00023_),
    .Q_N(_05643_),
    .Q(\uart0.txdiv[2] ));
 sg13g2_dfrbp_1 _13107_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00024_),
    .Q_N(_05642_),
    .Q(\uart0.txdiv[3] ));
 sg13g2_dfrbp_1 _13108_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00025_),
    .Q_N(_05641_),
    .Q(\uart0.txdiv[4] ));
 sg13g2_dfrbp_1 _13109_ (.CLK(net3916),
    .RESET_B(net3718),
    .D(_00026_),
    .Q_N(_05640_),
    .Q(\uart0.txdiv[5] ));
 sg13g2_tiehi _12449__18 (.L_HI(net18));
 sg13g2_tiehi _12448__19 (.L_HI(net19));
 sg13g2_tiehi _12447__20 (.L_HI(net20));
 sg13g2_tiehi _12446__21 (.L_HI(net21));
 sg13g2_tiehi _12445__22 (.L_HI(net22));
 sg13g2_tiehi _12444__23 (.L_HI(net23));
 sg13g2_tiehi _12443__24 (.L_HI(net24));
 sg13g2_tiehi _12442__25 (.L_HI(net25));
 sg13g2_tiehi _12441__26 (.L_HI(net26));
 sg13g2_tiehi _12440__27 (.L_HI(net27));
 sg13g2_tiehi _12439__28 (.L_HI(net28));
 sg13g2_tiehi _12438__29 (.L_HI(net29));
 sg13g2_tiehi _12437__30 (.L_HI(net30));
 sg13g2_tiehi _12436__31 (.L_HI(net31));
 sg13g2_tiehi _12435__32 (.L_HI(net32));
 sg13g2_tiehi _12434__33 (.L_HI(net33));
 sg13g2_tiehi _12433__34 (.L_HI(net34));
 sg13g2_tiehi _12432__35 (.L_HI(net35));
 sg13g2_tiehi _12431__36 (.L_HI(net36));
 sg13g2_tiehi _12430__37 (.L_HI(net37));
 sg13g2_tiehi _12429__38 (.L_HI(net38));
 sg13g2_tiehi _12428__39 (.L_HI(net39));
 sg13g2_tiehi _12427__40 (.L_HI(net40));
 sg13g2_tiehi _12426__41 (.L_HI(net41));
 sg13g2_tiehi _12425__42 (.L_HI(net42));
 sg13g2_tiehi _12424__43 (.L_HI(net43));
 sg13g2_tiehi _12423__44 (.L_HI(net44));
 sg13g2_tiehi _12422__45 (.L_HI(net45));
 sg13g2_tiehi _12421__46 (.L_HI(net46));
 sg13g2_tiehi _12420__47 (.L_HI(net47));
 sg13g2_tiehi _12419__48 (.L_HI(net48));
 sg13g2_tiehi _12418__49 (.L_HI(net49));
 sg13g2_tiehi _12417__50 (.L_HI(net50));
 sg13g2_tiehi _12416__51 (.L_HI(net51));
 sg13g2_tiehi _12415__52 (.L_HI(net52));
 sg13g2_tiehi _12414__53 (.L_HI(net53));
 sg13g2_tiehi _12413__54 (.L_HI(net54));
 sg13g2_tiehi _12412__55 (.L_HI(net55));
 sg13g2_tiehi _12411__56 (.L_HI(net56));
 sg13g2_tiehi _12410__57 (.L_HI(net57));
 sg13g2_tiehi _12409__58 (.L_HI(net58));
 sg13g2_tiehi _12408__59 (.L_HI(net59));
 sg13g2_tiehi _12407__60 (.L_HI(net60));
 sg13g2_tiehi _12406__61 (.L_HI(net61));
 sg13g2_tiehi _12405__62 (.L_HI(net62));
 sg13g2_tiehi _12404__63 (.L_HI(net63));
 sg13g2_tiehi _12403__64 (.L_HI(net64));
 sg13g2_tiehi _12402__65 (.L_HI(net65));
 sg13g2_tiehi _12401__66 (.L_HI(net66));
 sg13g2_tiehi _12400__67 (.L_HI(net67));
 sg13g2_tiehi _12399__68 (.L_HI(net68));
 sg13g2_tiehi _12398__69 (.L_HI(net69));
 sg13g2_tiehi _12397__70 (.L_HI(net70));
 sg13g2_tiehi _12396__71 (.L_HI(net71));
 sg13g2_tiehi _12395__72 (.L_HI(net72));
 sg13g2_tiehi _12394__73 (.L_HI(net73));
 sg13g2_tiehi _12393__74 (.L_HI(net74));
 sg13g2_tiehi _12392__75 (.L_HI(net75));
 sg13g2_tiehi _12391__76 (.L_HI(net76));
 sg13g2_tiehi _12390__77 (.L_HI(net77));
 sg13g2_tiehi _12389__78 (.L_HI(net78));
 sg13g2_tiehi _12388__79 (.L_HI(net79));
 sg13g2_tiehi _12387__80 (.L_HI(net80));
 sg13g2_tiehi _12386__81 (.L_HI(net81));
 sg13g2_tiehi _12385__82 (.L_HI(net82));
 sg13g2_tiehi _12384__83 (.L_HI(net83));
 sg13g2_tiehi _12383__84 (.L_HI(net84));
 sg13g2_tiehi _12382__85 (.L_HI(net85));
 sg13g2_tiehi _12381__86 (.L_HI(net86));
 sg13g2_tiehi _12380__87 (.L_HI(net87));
 sg13g2_tiehi _12379__88 (.L_HI(net88));
 sg13g2_tiehi _12378__89 (.L_HI(net89));
 sg13g2_tiehi _12377__90 (.L_HI(net90));
 sg13g2_tiehi _12376__91 (.L_HI(net91));
 sg13g2_tiehi _12375__92 (.L_HI(net92));
 sg13g2_tiehi _12374__93 (.L_HI(net93));
 sg13g2_tiehi _12373__94 (.L_HI(net94));
 sg13g2_tiehi _12372__95 (.L_HI(net95));
 sg13g2_tiehi _12371__96 (.L_HI(net96));
 sg13g2_tiehi _12370__97 (.L_HI(net97));
 sg13g2_tiehi _12369__98 (.L_HI(net98));
 sg13g2_tiehi _12368__99 (.L_HI(net99));
 sg13g2_tiehi _12367__100 (.L_HI(net100));
 sg13g2_tiehi _12366__101 (.L_HI(net101));
 sg13g2_tiehi _12365__102 (.L_HI(net102));
 sg13g2_tiehi _12364__103 (.L_HI(net103));
 sg13g2_tiehi _12363__104 (.L_HI(net104));
 sg13g2_tiehi _12362__105 (.L_HI(net105));
 sg13g2_tiehi _12361__106 (.L_HI(net106));
 sg13g2_tiehi _12360__107 (.L_HI(net107));
 sg13g2_tiehi _12359__108 (.L_HI(net108));
 sg13g2_tiehi _12358__109 (.L_HI(net109));
 sg13g2_tiehi _12357__110 (.L_HI(net110));
 sg13g2_tiehi _12356__111 (.L_HI(net111));
 sg13g2_tiehi _12355__112 (.L_HI(net112));
 sg13g2_tiehi _12354__113 (.L_HI(net113));
 sg13g2_tiehi _12353__114 (.L_HI(net114));
 sg13g2_tiehi _12352__115 (.L_HI(net115));
 sg13g2_tiehi _12351__116 (.L_HI(net116));
 sg13g2_tiehi _12350__117 (.L_HI(net117));
 sg13g2_tiehi _12349__118 (.L_HI(net118));
 sg13g2_tiehi _12348__119 (.L_HI(net119));
 sg13g2_tiehi _12347__120 (.L_HI(net120));
 sg13g2_tiehi _12346__121 (.L_HI(net121));
 sg13g2_tiehi _12345__122 (.L_HI(net122));
 sg13g2_tiehi _12344__123 (.L_HI(net123));
 sg13g2_tiehi _12343__124 (.L_HI(net124));
 sg13g2_tiehi _12342__125 (.L_HI(net125));
 sg13g2_tiehi _12341__126 (.L_HI(net126));
 sg13g2_tiehi _12340__127 (.L_HI(net127));
 sg13g2_tiehi _12339__128 (.L_HI(net128));
 sg13g2_tiehi _12338__129 (.L_HI(net129));
 sg13g2_tiehi _12337__130 (.L_HI(net130));
 sg13g2_tiehi _12336__131 (.L_HI(net131));
 sg13g2_tiehi _12335__132 (.L_HI(net132));
 sg13g2_tiehi _12334__133 (.L_HI(net133));
 sg13g2_tiehi _12333__134 (.L_HI(net134));
 sg13g2_tiehi _12332__135 (.L_HI(net135));
 sg13g2_tiehi _12331__136 (.L_HI(net136));
 sg13g2_tiehi _12330__137 (.L_HI(net137));
 sg13g2_tiehi _12329__138 (.L_HI(net138));
 sg13g2_tiehi _12328__139 (.L_HI(net139));
 sg13g2_tiehi _12327__140 (.L_HI(net140));
 sg13g2_tiehi _12326__141 (.L_HI(net141));
 sg13g2_tiehi _12325__142 (.L_HI(net142));
 sg13g2_tiehi _12324__143 (.L_HI(net143));
 sg13g2_tiehi _12323__144 (.L_HI(net144));
 sg13g2_tiehi _12322__145 (.L_HI(net145));
 sg13g2_tiehi _12321__146 (.L_HI(net146));
 sg13g2_tiehi _12320__147 (.L_HI(net147));
 sg13g2_tiehi _12319__148 (.L_HI(net148));
 sg13g2_tiehi _12318__149 (.L_HI(net149));
 sg13g2_tiehi _12317__150 (.L_HI(net150));
 sg13g2_tiehi _12316__151 (.L_HI(net151));
 sg13g2_tiehi _12315__152 (.L_HI(net152));
 sg13g2_tiehi _12314__153 (.L_HI(net153));
 sg13g2_tiehi _12313__154 (.L_HI(net154));
 sg13g2_tiehi _12312__155 (.L_HI(net155));
 sg13g2_tiehi _12311__156 (.L_HI(net156));
 sg13g2_tiehi _12310__157 (.L_HI(net157));
 sg13g2_tiehi _12309__158 (.L_HI(net158));
 sg13g2_tiehi _12308__159 (.L_HI(net159));
 sg13g2_tiehi _12307__160 (.L_HI(net160));
 sg13g2_tiehi _12306__161 (.L_HI(net161));
 sg13g2_tiehi _12305__162 (.L_HI(net162));
 sg13g2_tiehi _12304__163 (.L_HI(net163));
 sg13g2_tiehi _12303__164 (.L_HI(net164));
 sg13g2_tiehi _12302__165 (.L_HI(net165));
 sg13g2_tiehi _12301__166 (.L_HI(net166));
 sg13g2_tiehi _12300__167 (.L_HI(net167));
 sg13g2_tiehi _12299__168 (.L_HI(net168));
 sg13g2_tiehi _12298__169 (.L_HI(net169));
 sg13g2_tiehi _12297__170 (.L_HI(net170));
 sg13g2_tiehi _12296__171 (.L_HI(net171));
 sg13g2_tiehi _12295__172 (.L_HI(net172));
 sg13g2_tiehi _12294__173 (.L_HI(net173));
 sg13g2_tiehi _12293__174 (.L_HI(net174));
 sg13g2_tiehi _12292__175 (.L_HI(net175));
 sg13g2_tiehi _12291__176 (.L_HI(net176));
 sg13g2_tiehi _12290__177 (.L_HI(net177));
 sg13g2_tiehi _12289__178 (.L_HI(net178));
 sg13g2_tiehi _12288__179 (.L_HI(net179));
 sg13g2_tiehi _12287__180 (.L_HI(net180));
 sg13g2_tiehi _12286__181 (.L_HI(net181));
 sg13g2_tiehi _12285__182 (.L_HI(net182));
 sg13g2_tiehi _12284__183 (.L_HI(net183));
 sg13g2_tiehi _12283__184 (.L_HI(net184));
 sg13g2_tiehi _12282__185 (.L_HI(net185));
 sg13g2_tiehi _12281__186 (.L_HI(net186));
 sg13g2_tiehi _12280__187 (.L_HI(net187));
 sg13g2_tiehi _12279__188 (.L_HI(net188));
 sg13g2_tiehi _12278__189 (.L_HI(net189));
 sg13g2_tiehi _12277__190 (.L_HI(net190));
 sg13g2_tiehi _12276__191 (.L_HI(net191));
 sg13g2_tiehi _12275__192 (.L_HI(net192));
 sg13g2_tiehi _12274__193 (.L_HI(net193));
 sg13g2_tiehi _12273__194 (.L_HI(net194));
 sg13g2_tiehi _12272__195 (.L_HI(net195));
 sg13g2_tiehi _12271__196 (.L_HI(net196));
 sg13g2_tiehi _12270__197 (.L_HI(net197));
 sg13g2_tiehi _12269__198 (.L_HI(net198));
 sg13g2_tiehi _12268__199 (.L_HI(net199));
 sg13g2_tiehi _12267__200 (.L_HI(net200));
 sg13g2_tiehi _12266__201 (.L_HI(net201));
 sg13g2_tiehi _12265__202 (.L_HI(net202));
 sg13g2_tiehi _12264__203 (.L_HI(net203));
 sg13g2_tiehi _12263__204 (.L_HI(net204));
 sg13g2_tiehi _12262__205 (.L_HI(net205));
 sg13g2_tiehi _12261__206 (.L_HI(net206));
 sg13g2_tiehi _12260__207 (.L_HI(net207));
 sg13g2_tiehi _12259__208 (.L_HI(net208));
 sg13g2_tiehi _12258__209 (.L_HI(net209));
 sg13g2_tiehi _12257__210 (.L_HI(net210));
 sg13g2_tiehi _12256__211 (.L_HI(net211));
 sg13g2_tiehi _12255__212 (.L_HI(net212));
 sg13g2_tiehi _12254__213 (.L_HI(net213));
 sg13g2_tiehi _12253__214 (.L_HI(net214));
 sg13g2_tiehi _12252__215 (.L_HI(net215));
 sg13g2_tiehi _12251__216 (.L_HI(net216));
 sg13g2_tiehi _12250__217 (.L_HI(net217));
 sg13g2_tiehi _12249__218 (.L_HI(net218));
 sg13g2_tiehi _12248__219 (.L_HI(net219));
 sg13g2_tiehi _12247__220 (.L_HI(net220));
 sg13g2_tiehi _12246__221 (.L_HI(net221));
 sg13g2_tiehi _12245__222 (.L_HI(net222));
 sg13g2_tiehi _12244__223 (.L_HI(net223));
 sg13g2_tiehi _12243__224 (.L_HI(net224));
 sg13g2_tiehi _12242__225 (.L_HI(net225));
 sg13g2_tiehi _12241__226 (.L_HI(net226));
 sg13g2_tiehi _12240__227 (.L_HI(net227));
 sg13g2_tiehi _12239__228 (.L_HI(net228));
 sg13g2_tiehi _12238__229 (.L_HI(net229));
 sg13g2_tiehi _12237__230 (.L_HI(net230));
 sg13g2_tiehi _12236__231 (.L_HI(net231));
 sg13g2_tiehi _12235__232 (.L_HI(net232));
 sg13g2_tiehi _12234__233 (.L_HI(net233));
 sg13g2_tiehi _12233__234 (.L_HI(net234));
 sg13g2_tiehi _12232__235 (.L_HI(net235));
 sg13g2_tiehi _12231__236 (.L_HI(net236));
 sg13g2_tiehi _12230__237 (.L_HI(net237));
 sg13g2_tiehi _12229__238 (.L_HI(net238));
 sg13g2_tiehi _12228__239 (.L_HI(net239));
 sg13g2_tiehi _12227__240 (.L_HI(net240));
 sg13g2_tiehi _12226__241 (.L_HI(net241));
 sg13g2_tiehi _12225__242 (.L_HI(net242));
 sg13g2_tiehi _12224__243 (.L_HI(net243));
 sg13g2_tiehi _12223__244 (.L_HI(net244));
 sg13g2_tiehi _12222__245 (.L_HI(net245));
 sg13g2_tiehi _12221__246 (.L_HI(net246));
 sg13g2_tiehi _12220__247 (.L_HI(net247));
 sg13g2_tiehi _12219__248 (.L_HI(net248));
 sg13g2_tiehi _12218__249 (.L_HI(net249));
 sg13g2_tiehi _12217__250 (.L_HI(net250));
 sg13g2_tiehi _12216__251 (.L_HI(net251));
 sg13g2_tiehi _12215__252 (.L_HI(net252));
 sg13g2_tiehi _12214__253 (.L_HI(net253));
 sg13g2_tiehi _12213__254 (.L_HI(net254));
 sg13g2_tiehi _12212__255 (.L_HI(net255));
 sg13g2_tiehi _12211__256 (.L_HI(net256));
 sg13g2_tiehi _12210__257 (.L_HI(net257));
 sg13g2_tiehi _12209__258 (.L_HI(net258));
 sg13g2_tiehi _12208__259 (.L_HI(net259));
 sg13g2_tiehi _12207__260 (.L_HI(net260));
 sg13g2_tiehi _12206__261 (.L_HI(net261));
 sg13g2_tiehi _12205__262 (.L_HI(net262));
 sg13g2_tiehi _12204__263 (.L_HI(net263));
 sg13g2_tiehi _12203__264 (.L_HI(net264));
 sg13g2_tiehi _12202__265 (.L_HI(net265));
 sg13g2_tiehi _12201__266 (.L_HI(net266));
 sg13g2_tiehi _12200__267 (.L_HI(net267));
 sg13g2_tiehi _12199__268 (.L_HI(net268));
 sg13g2_tiehi _12198__269 (.L_HI(net269));
 sg13g2_tiehi _12197__270 (.L_HI(net270));
 sg13g2_tiehi _12196__271 (.L_HI(net271));
 sg13g2_tiehi _12195__272 (.L_HI(net272));
 sg13g2_tiehi _12194__273 (.L_HI(net273));
 sg13g2_tiehi _12193__274 (.L_HI(net274));
 sg13g2_tiehi _12192__275 (.L_HI(net275));
 sg13g2_tiehi _12191__276 (.L_HI(net276));
 sg13g2_tiehi _12190__277 (.L_HI(net277));
 sg13g2_tiehi _12189__278 (.L_HI(net278));
 sg13g2_tiehi _12188__279 (.L_HI(net279));
 sg13g2_tiehi _12187__280 (.L_HI(net280));
 sg13g2_tiehi _12186__281 (.L_HI(net281));
 sg13g2_tiehi _12185__282 (.L_HI(net282));
 sg13g2_tiehi _12184__283 (.L_HI(net283));
 sg13g2_tiehi _12183__284 (.L_HI(net284));
 sg13g2_tiehi _12182__285 (.L_HI(net285));
 sg13g2_tiehi _12181__286 (.L_HI(net286));
 sg13g2_tiehi _12180__287 (.L_HI(net287));
 sg13g2_tiehi _12179__288 (.L_HI(net288));
 sg13g2_tiehi _12178__289 (.L_HI(net289));
 sg13g2_tiehi _12177__290 (.L_HI(net290));
 sg13g2_tiehi _12176__291 (.L_HI(net291));
 sg13g2_tiehi _12175__292 (.L_HI(net292));
 sg13g2_tiehi _12174__293 (.L_HI(net293));
 sg13g2_tiehi _12173__294 (.L_HI(net294));
 sg13g2_tiehi _12172__295 (.L_HI(net295));
 sg13g2_tiehi _12171__296 (.L_HI(net296));
 sg13g2_tiehi _12170__297 (.L_HI(net297));
 sg13g2_tiehi _12169__298 (.L_HI(net298));
 sg13g2_tiehi _12168__299 (.L_HI(net299));
 sg13g2_tiehi _12167__300 (.L_HI(net300));
 sg13g2_tiehi _12166__301 (.L_HI(net301));
 sg13g2_tiehi _12165__302 (.L_HI(net302));
 sg13g2_tiehi _12164__303 (.L_HI(net303));
 sg13g2_tiehi _12163__304 (.L_HI(net304));
 sg13g2_tiehi _12162__305 (.L_HI(net305));
 sg13g2_tiehi _12161__306 (.L_HI(net306));
 sg13g2_tiehi _12160__307 (.L_HI(net307));
 sg13g2_tiehi _12159__308 (.L_HI(net308));
 sg13g2_tiehi _12158__309 (.L_HI(net309));
 sg13g2_tiehi _12157__310 (.L_HI(net310));
 sg13g2_tiehi _12156__311 (.L_HI(net311));
 sg13g2_tiehi _12155__312 (.L_HI(net312));
 sg13g2_tiehi _12154__313 (.L_HI(net313));
 sg13g2_tiehi _12153__314 (.L_HI(net314));
 sg13g2_tiehi _12152__315 (.L_HI(net315));
 sg13g2_tiehi _12151__316 (.L_HI(net316));
 sg13g2_tiehi _12150__317 (.L_HI(net317));
 sg13g2_tiehi _12149__318 (.L_HI(net318));
 sg13g2_tiehi _12148__319 (.L_HI(net319));
 sg13g2_tiehi _12147__320 (.L_HI(net320));
 sg13g2_tiehi _12146__321 (.L_HI(net321));
 sg13g2_tiehi _12145__322 (.L_HI(net322));
 sg13g2_tiehi _12144__323 (.L_HI(net323));
 sg13g2_tiehi _12143__324 (.L_HI(net324));
 sg13g2_tiehi _12142__325 (.L_HI(net325));
 sg13g2_tiehi _12141__326 (.L_HI(net326));
 sg13g2_tiehi _12140__327 (.L_HI(net327));
 sg13g2_tiehi _12889__328 (.L_HI(net328));
 sg13g2_tiehi _12888__329 (.L_HI(net329));
 sg13g2_tiehi _12887__330 (.L_HI(net330));
 sg13g2_tiehi _12886__331 (.L_HI(net331));
 sg13g2_tiehi _12885__332 (.L_HI(net332));
 sg13g2_tiehi _12884__333 (.L_HI(net333));
 sg13g2_tiehi _12883__334 (.L_HI(net334));
 sg13g2_tiehi _12882__335 (.L_HI(net335));
 sg13g2_tiehi _12881__336 (.L_HI(net336));
 sg13g2_tiehi _12880__337 (.L_HI(net337));
 sg13g2_tiehi _12879__338 (.L_HI(net338));
 sg13g2_tiehi _12878__339 (.L_HI(net339));
 sg13g2_tiehi _12877__340 (.L_HI(net340));
 sg13g2_tiehi _12876__341 (.L_HI(net341));
 sg13g2_tiehi _12875__342 (.L_HI(net342));
 sg13g2_tiehi _12874__343 (.L_HI(net343));
 sg13g2_tiehi _12873__344 (.L_HI(net344));
 sg13g2_tiehi _12872__345 (.L_HI(net345));
 sg13g2_tiehi _12871__346 (.L_HI(net346));
 sg13g2_tiehi _12870__347 (.L_HI(net347));
 sg13g2_tiehi _12869__348 (.L_HI(net348));
 sg13g2_tiehi _12868__349 (.L_HI(net349));
 sg13g2_tiehi _12867__350 (.L_HI(net350));
 sg13g2_tiehi _12866__351 (.L_HI(net351));
 sg13g2_tiehi _12865__352 (.L_HI(net352));
 sg13g2_tiehi _12864__353 (.L_HI(net353));
 sg13g2_tiehi _12863__354 (.L_HI(net354));
 sg13g2_tiehi _12862__355 (.L_HI(net355));
 sg13g2_tiehi _12861__356 (.L_HI(net356));
 sg13g2_tiehi _12860__357 (.L_HI(net357));
 sg13g2_tiehi _12859__358 (.L_HI(net358));
 sg13g2_tiehi _12858__359 (.L_HI(net359));
 sg13g2_tiehi _12857__360 (.L_HI(net360));
 sg13g2_tiehi _12856__361 (.L_HI(net361));
 sg13g2_tiehi _12855__362 (.L_HI(net362));
 sg13g2_tiehi _12854__363 (.L_HI(net363));
 sg13g2_tiehi _12853__364 (.L_HI(net364));
 sg13g2_tiehi _12852__365 (.L_HI(net365));
 sg13g2_tiehi _12851__366 (.L_HI(net366));
 sg13g2_tiehi _12850__367 (.L_HI(net367));
 sg13g2_tiehi _12849__368 (.L_HI(net368));
 sg13g2_tiehi _12848__369 (.L_HI(net369));
 sg13g2_tiehi _12847__370 (.L_HI(net370));
 sg13g2_tiehi _12846__371 (.L_HI(net371));
 sg13g2_tiehi _12845__372 (.L_HI(net372));
 sg13g2_tiehi _12844__373 (.L_HI(net373));
 sg13g2_tiehi _12843__374 (.L_HI(net374));
 sg13g2_tiehi _12842__375 (.L_HI(net375));
 sg13g2_tiehi _12841__376 (.L_HI(net376));
 sg13g2_tiehi _12840__377 (.L_HI(net377));
 sg13g2_tiehi _12839__378 (.L_HI(net378));
 sg13g2_tiehi _12838__379 (.L_HI(net379));
 sg13g2_tiehi _12837__380 (.L_HI(net380));
 sg13g2_tiehi _12836__381 (.L_HI(net381));
 sg13g2_tiehi _12835__382 (.L_HI(net382));
 sg13g2_tiehi _13096__383 (.L_HI(net383));
 sg13g2_tiehi _12834__384 (.L_HI(net384));
 sg13g2_tiehi _12833__385 (.L_HI(net385));
 sg13g2_tiehi _12832__386 (.L_HI(net386));
 sg13g2_tiehi _13095__387 (.L_HI(net387));
 sg13g2_tiehi _12831__388 (.L_HI(net388));
 sg13g2_tiehi _12830__389 (.L_HI(net389));
 sg13g2_tiehi _12829__390 (.L_HI(net390));
 sg13g2_tiehi _13094__391 (.L_HI(net391));
 sg13g2_tiehi _12828__392 (.L_HI(net392));
 sg13g2_tiehi _13103__393 (.L_HI(net393));
 sg13g2_tiehi _12827__394 (.L_HI(net394));
 sg13g2_tiehi _13093__395 (.L_HI(net395));
 sg13g2_tiehi _12826__396 (.L_HI(net396));
 sg13g2_tiehi _12825__397 (.L_HI(net397));
 sg13g2_tiehi _12824__398 (.L_HI(net398));
 sg13g2_tiehi _13092__399 (.L_HI(net399));
 sg13g2_tiehi _12823__400 (.L_HI(net400));
 sg13g2_tiehi _13102__401 (.L_HI(net401));
 sg13g2_tiehi _12822__402 (.L_HI(net402));
 sg13g2_tiehi _12821__403 (.L_HI(net403));
 sg13g2_tiehi _13091__404 (.L_HI(net404));
 sg13g2_tiehi _12820__405 (.L_HI(net405));
 sg13g2_tiehi _12819__406 (.L_HI(net406));
 sg13g2_tiehi _13090__407 (.L_HI(net407));
 sg13g2_tiehi _12818__408 (.L_HI(net408));
 sg13g2_tiehi _12817__409 (.L_HI(net409));
 sg13g2_tiehi _13101__410 (.L_HI(net410));
 sg13g2_tiehi _12816__411 (.L_HI(net411));
 sg13g2_tiehi _13089__412 (.L_HI(net412));
 sg13g2_tiehi _12815__413 (.L_HI(net413));
 sg13g2_tiehi _12814__414 (.L_HI(net414));
 sg13g2_tiehi _12813__415 (.L_HI(net415));
 sg13g2_tiehi _13088__416 (.L_HI(net416));
 sg13g2_tiehi _12812__417 (.L_HI(net417));
 sg13g2_tiehi _12139__418 (.L_HI(net418));
 sg13g2_tiehi _12811__419 (.L_HI(net419));
 sg13g2_tiehi _12810__420 (.L_HI(net420));
 sg13g2_tiehi _12809__421 (.L_HI(net421));
 sg13g2_tiehi _12808__422 (.L_HI(net422));
 sg13g2_tiehi _12807__423 (.L_HI(net423));
 sg13g2_tiehi _12806__424 (.L_HI(net424));
 sg13g2_tiehi _12805__425 (.L_HI(net425));
 sg13g2_tiehi _12804__426 (.L_HI(net426));
 sg13g2_tiehi _12803__427 (.L_HI(net427));
 sg13g2_tiehi _12802__428 (.L_HI(net428));
 sg13g2_tiehi _12801__429 (.L_HI(net429));
 sg13g2_tiehi _13068__430 (.L_HI(net430));
 sg13g2_tiehi _12800__431 (.L_HI(net431));
 sg13g2_tiehi _13067__432 (.L_HI(net432));
 sg13g2_tiehi _12799__433 (.L_HI(net433));
 sg13g2_tiehi _13066__434 (.L_HI(net434));
 sg13g2_tiehi _12798__435 (.L_HI(net435));
 sg13g2_tiehi _13065__436 (.L_HI(net436));
 sg13g2_tiehi _12797__437 (.L_HI(net437));
 sg13g2_tiehi _13064__438 (.L_HI(net438));
 sg13g2_tiehi _12796__439 (.L_HI(net439));
 sg13g2_tiehi _13063__440 (.L_HI(net440));
 sg13g2_tiehi _12795__441 (.L_HI(net441));
 sg13g2_tiehi _13062__442 (.L_HI(net442));
 sg13g2_tiehi _12794__443 (.L_HI(net443));
 sg13g2_tiehi _13061__444 (.L_HI(net444));
 sg13g2_tiehi _12793__445 (.L_HI(net445));
 sg13g2_tiehi _13060__446 (.L_HI(net446));
 sg13g2_tiehi _12792__447 (.L_HI(net447));
 sg13g2_tiehi _13059__448 (.L_HI(net448));
 sg13g2_tiehi _12791__449 (.L_HI(net449));
 sg13g2_tiehi _13058__450 (.L_HI(net450));
 sg13g2_tiehi _12790__451 (.L_HI(net451));
 sg13g2_tiehi _13057__452 (.L_HI(net452));
 sg13g2_tiehi _12789__453 (.L_HI(net453));
 sg13g2_tiehi _13056__454 (.L_HI(net454));
 sg13g2_tiehi _12788__455 (.L_HI(net455));
 sg13g2_tiehi _13055__456 (.L_HI(net456));
 sg13g2_tiehi _12787__457 (.L_HI(net457));
 sg13g2_tiehi _13054__458 (.L_HI(net458));
 sg13g2_tiehi _12786__459 (.L_HI(net459));
 sg13g2_tiehi _13053__460 (.L_HI(net460));
 sg13g2_tiehi _12785__461 (.L_HI(net461));
 sg13g2_tiehi _13052__462 (.L_HI(net462));
 sg13g2_tiehi _12784__463 (.L_HI(net463));
 sg13g2_tiehi _13051__464 (.L_HI(net464));
 sg13g2_tiehi _12783__465 (.L_HI(net465));
 sg13g2_tiehi _13050__466 (.L_HI(net466));
 sg13g2_tiehi _12782__467 (.L_HI(net467));
 sg13g2_tiehi _13049__468 (.L_HI(net468));
 sg13g2_tiehi _12781__469 (.L_HI(net469));
 sg13g2_tiehi _13048__470 (.L_HI(net470));
 sg13g2_tiehi _13047__471 (.L_HI(net471));
 sg13g2_tiehi _12780__472 (.L_HI(net472));
 sg13g2_tiehi _13046__473 (.L_HI(net473));
 sg13g2_tiehi _13045__474 (.L_HI(net474));
 sg13g2_tiehi _12779__475 (.L_HI(net475));
 sg13g2_tiehi _13044__476 (.L_HI(net476));
 sg13g2_tiehi _13043__477 (.L_HI(net477));
 sg13g2_tiehi _12778__478 (.L_HI(net478));
 sg13g2_tiehi _13042__479 (.L_HI(net479));
 sg13g2_tiehi _13041__480 (.L_HI(net480));
 sg13g2_tiehi _12637__481 (.L_HI(net481));
 sg13g2_tiehi _12777__482 (.L_HI(net482));
 sg13g2_tiehi _13040__483 (.L_HI(net483));
 sg13g2_tiehi _13039__484 (.L_HI(net484));
 sg13g2_tiehi _12776__485 (.L_HI(net485));
 sg13g2_tiehi _12775__486 (.L_HI(net486));
 sg13g2_tiehi _12774__487 (.L_HI(net487));
 sg13g2_tiehi _12773__488 (.L_HI(net488));
 sg13g2_tiehi _12772__489 (.L_HI(net489));
 sg13g2_tiehi _12771__490 (.L_HI(net490));
 sg13g2_tiehi _12770__491 (.L_HI(net491));
 sg13g2_tiehi _12769__492 (.L_HI(net492));
 sg13g2_tiehi _12768__493 (.L_HI(net493));
 sg13g2_tiehi _12767__494 (.L_HI(net494));
 sg13g2_tiehi _12766__495 (.L_HI(net495));
 sg13g2_tiehi _12765__496 (.L_HI(net496));
 sg13g2_tiehi _12764__497 (.L_HI(net497));
 sg13g2_tiehi _12763__498 (.L_HI(net498));
 sg13g2_tiehi _12762__499 (.L_HI(net499));
 sg13g2_tiehi _12761__500 (.L_HI(net500));
 sg13g2_tiehi _12976__501 (.L_HI(net501));
 sg13g2_tiehi _12942__502 (.L_HI(net502));
 sg13g2_tiehi _12760__503 (.L_HI(net503));
 sg13g2_tiehi _12941__504 (.L_HI(net504));
 sg13g2_tiehi _12940__505 (.L_HI(net505));
 sg13g2_tiehi _12759__506 (.L_HI(net506));
 sg13g2_tiehi _12939__507 (.L_HI(net507));
 sg13g2_tiehi _12938__508 (.L_HI(net508));
 sg13g2_tiehi _12758__509 (.L_HI(net509));
 sg13g2_tiehi _12937__510 (.L_HI(net510));
 sg13g2_tiehi _12936__511 (.L_HI(net511));
 sg13g2_tiehi _12757__512 (.L_HI(net512));
 sg13g2_tiehi _12756__513 (.L_HI(net513));
 sg13g2_tiehi _12934__514 (.L_HI(net514));
 sg13g2_tiehi _12755__515 (.L_HI(net515));
 sg13g2_tiehi _12933__516 (.L_HI(net516));
 sg13g2_tiehi _12932__517 (.L_HI(net517));
 sg13g2_tiehi _12754__518 (.L_HI(net518));
 sg13g2_tiehi _12931__519 (.L_HI(net519));
 sg13g2_tiehi _12930__520 (.L_HI(net520));
 sg13g2_tiehi _12753__521 (.L_HI(net521));
 sg13g2_tiehi _12929__522 (.L_HI(net522));
 sg13g2_tiehi _12928__523 (.L_HI(net523));
 sg13g2_tiehi _12752__524 (.L_HI(net524));
 sg13g2_tiehi _12927__525 (.L_HI(net525));
 sg13g2_tiehi _12926__526 (.L_HI(net526));
 sg13g2_tiehi _12751__527 (.L_HI(net527));
 sg13g2_tiehi _12925__528 (.L_HI(net528));
 sg13g2_tiehi _12924__529 (.L_HI(net529));
 sg13g2_tiehi _12750__530 (.L_HI(net530));
 sg13g2_tiehi _12923__531 (.L_HI(net531));
 sg13g2_tiehi _12922__532 (.L_HI(net532));
 sg13g2_tiehi _12749__533 (.L_HI(net533));
 sg13g2_tiehi _12921__534 (.L_HI(net534));
 sg13g2_tiehi _12748__535 (.L_HI(net535));
 sg13g2_tiehi _12920__536 (.L_HI(net536));
 sg13g2_tiehi _12919__537 (.L_HI(net537));
 sg13g2_tiehi _12918__538 (.L_HI(net538));
 sg13g2_tiehi _12743__539 (.L_HI(net539));
 sg13g2_tiehi _12738__540 (.L_HI(net540));
 sg13g2_tiehi _12737__541 (.L_HI(net541));
 sg13g2_tiehi _12736__542 (.L_HI(net542));
 sg13g2_tiehi _12641__543 (.L_HI(net543));
 sg13g2_tiehi _12735__544 (.L_HI(net544));
 sg13g2_tiehi _12734__545 (.L_HI(net545));
 sg13g2_tiehi _12733__546 (.L_HI(net546));
 sg13g2_tiehi _12732__547 (.L_HI(net547));
 sg13g2_tiehi _12731__548 (.L_HI(net548));
 sg13g2_tiehi _12730__549 (.L_HI(net549));
 sg13g2_tiehi _12729__550 (.L_HI(net550));
 sg13g2_tiehi _12728__551 (.L_HI(net551));
 sg13g2_tiehi _12727__552 (.L_HI(net552));
 sg13g2_tiehi _12726__553 (.L_HI(net553));
 sg13g2_tiehi _12725__554 (.L_HI(net554));
 sg13g2_tiehi _12724__555 (.L_HI(net555));
 sg13g2_tiehi _12723__556 (.L_HI(net556));
 sg13g2_tiehi _12722__557 (.L_HI(net557));
 sg13g2_tiehi _12721__558 (.L_HI(net558));
 sg13g2_tiehi _12720__559 (.L_HI(net559));
 sg13g2_tiehi _12719__560 (.L_HI(net560));
 sg13g2_tiehi _12718__561 (.L_HI(net561));
 sg13g2_tiehi _12717__562 (.L_HI(net562));
 sg13g2_tiehi _12716__563 (.L_HI(net563));
 sg13g2_tiehi _12715__564 (.L_HI(net564));
 sg13g2_tiehi _12714__565 (.L_HI(net565));
 sg13g2_tiehi _12713__566 (.L_HI(net566));
 sg13g2_tiehi _12712__567 (.L_HI(net567));
 sg13g2_tiehi _12711__568 (.L_HI(net568));
 sg13g2_tiehi _12710__569 (.L_HI(net569));
 sg13g2_tiehi _12709__570 (.L_HI(net570));
 sg13g2_tiehi _12708__571 (.L_HI(net571));
 sg13g2_tiehi _12707__572 (.L_HI(net572));
 sg13g2_tiehi _12706__573 (.L_HI(net573));
 sg13g2_tiehi _12705__574 (.L_HI(net574));
 sg13g2_tiehi _12704__575 (.L_HI(net575));
 sg13g2_tiehi _12703__576 (.L_HI(net576));
 sg13g2_tiehi _12702__577 (.L_HI(net577));
 sg13g2_tiehi _12701__578 (.L_HI(net578));
 sg13g2_tiehi _12700__579 (.L_HI(net579));
 sg13g2_tiehi _12699__580 (.L_HI(net580));
 sg13g2_tiehi _12698__581 (.L_HI(net581));
 sg13g2_tiehi _12697__582 (.L_HI(net582));
 sg13g2_tiehi _12696__583 (.L_HI(net583));
 sg13g2_tiehi _12695__584 (.L_HI(net584));
 sg13g2_tiehi _12694__585 (.L_HI(net585));
 sg13g2_tiehi _12693__586 (.L_HI(net586));
 sg13g2_tiehi _12692__587 (.L_HI(net587));
 sg13g2_tiehi _12691__588 (.L_HI(net588));
 sg13g2_tiehi _12690__589 (.L_HI(net589));
 sg13g2_tiehi _12689__590 (.L_HI(net590));
 sg13g2_tiehi _12688__591 (.L_HI(net591));
 sg13g2_tiehi _12687__592 (.L_HI(net592));
 sg13g2_tiehi _12686__593 (.L_HI(net593));
 sg13g2_tiehi _12685__594 (.L_HI(net594));
 sg13g2_tiehi _12684__595 (.L_HI(net595));
 sg13g2_tiehi _12683__596 (.L_HI(net596));
 sg13g2_tiehi _12682__597 (.L_HI(net597));
 sg13g2_tiehi _12681__598 (.L_HI(net598));
 sg13g2_tiehi _12680__599 (.L_HI(net599));
 sg13g2_tiehi _12679__600 (.L_HI(net600));
 sg13g2_tiehi _12678__601 (.L_HI(net601));
 sg13g2_tiehi _12677__602 (.L_HI(net602));
 sg13g2_tiehi _12676__603 (.L_HI(net603));
 sg13g2_tiehi _12675__604 (.L_HI(net604));
 sg13g2_tiehi _12674__605 (.L_HI(net605));
 sg13g2_tiehi _12673__606 (.L_HI(net606));
 sg13g2_tiehi _12672__607 (.L_HI(net607));
 sg13g2_tiehi _12671__608 (.L_HI(net608));
 sg13g2_tiehi _12670__609 (.L_HI(net609));
 sg13g2_tiehi _12669__610 (.L_HI(net610));
 sg13g2_tiehi _12668__611 (.L_HI(net611));
 sg13g2_tiehi _12667__612 (.L_HI(net612));
 sg13g2_tiehi _12666__613 (.L_HI(net613));
 sg13g2_tiehi _12665__614 (.L_HI(net614));
 sg13g2_tiehi _12664__615 (.L_HI(net615));
 sg13g2_tiehi _12663__616 (.L_HI(net616));
 sg13g2_tiehi _12662__617 (.L_HI(net617));
 sg13g2_tiehi _12661__618 (.L_HI(net618));
 sg13g2_tiehi _12660__619 (.L_HI(net619));
 sg13g2_tiehi _12659__620 (.L_HI(net620));
 sg13g2_tiehi _12658__621 (.L_HI(net621));
 sg13g2_tiehi _12657__622 (.L_HI(net622));
 sg13g2_tiehi _12656__623 (.L_HI(net623));
 sg13g2_tiehi _12655__624 (.L_HI(net624));
 sg13g2_tiehi _12654__625 (.L_HI(net625));
 sg13g2_tiehi _12653__626 (.L_HI(net626));
 sg13g2_tiehi _12652__627 (.L_HI(net627));
 sg13g2_tiehi _12651__628 (.L_HI(net628));
 sg13g2_tiehi _12650__629 (.L_HI(net629));
 sg13g2_tiehi _12649__630 (.L_HI(net630));
 sg13g2_tiehi _12648__631 (.L_HI(net631));
 sg13g2_tiehi _12647__632 (.L_HI(net632));
 sg13g2_tiehi _12646__633 (.L_HI(net633));
 sg13g2_tiehi _12645__634 (.L_HI(net634));
 sg13g2_tiehi _12644__635 (.L_HI(net635));
 sg13g2_tiehi _12643__636 (.L_HI(net636));
 sg13g2_tiehi _12636__637 (.L_HI(net637));
 sg13g2_tiehi _12635__638 (.L_HI(net638));
 sg13g2_tiehi _12634__639 (.L_HI(net639));
 sg13g2_tiehi _12633__640 (.L_HI(net640));
 sg13g2_tiehi _12632__641 (.L_HI(net641));
 sg13g2_tiehi _12631__642 (.L_HI(net642));
 sg13g2_tiehi _12630__643 (.L_HI(net643));
 sg13g2_tiehi _12629__644 (.L_HI(net644));
 sg13g2_tiehi _12628__645 (.L_HI(net645));
 sg13g2_tiehi _12627__646 (.L_HI(net646));
 sg13g2_tiehi _12626__647 (.L_HI(net647));
 sg13g2_tiehi _12625__648 (.L_HI(net648));
 sg13g2_tiehi _12624__649 (.L_HI(net649));
 sg13g2_tiehi _12623__650 (.L_HI(net650));
 sg13g2_tiehi _12622__651 (.L_HI(net651));
 sg13g2_tiehi _12620__652 (.L_HI(net652));
 sg13g2_tiehi _12619__653 (.L_HI(net653));
 sg13g2_tiehi _12618__654 (.L_HI(net654));
 sg13g2_tiehi _12617__655 (.L_HI(net655));
 sg13g2_tiehi _12616__656 (.L_HI(net656));
 sg13g2_tiehi _12615__657 (.L_HI(net657));
 sg13g2_tiehi _12614__658 (.L_HI(net658));
 sg13g2_tiehi _12613__659 (.L_HI(net659));
 sg13g2_tiehi _12612__660 (.L_HI(net660));
 sg13g2_tiehi _12611__661 (.L_HI(net661));
 sg13g2_tiehi _12610__662 (.L_HI(net662));
 sg13g2_tiehi _12609__663 (.L_HI(net663));
 sg13g2_tiehi _12608__664 (.L_HI(net664));
 sg13g2_tiehi _12607__665 (.L_HI(net665));
 sg13g2_tiehi _12606__666 (.L_HI(net666));
 sg13g2_tiehi _12605__667 (.L_HI(net667));
 sg13g2_tiehi _12604__668 (.L_HI(net668));
 sg13g2_tiehi _12603__669 (.L_HI(net669));
 sg13g2_tiehi _12602__670 (.L_HI(net670));
 sg13g2_tiehi _12601__671 (.L_HI(net671));
 sg13g2_tiehi _12600__672 (.L_HI(net672));
 sg13g2_tiehi _12599__673 (.L_HI(net673));
 sg13g2_tiehi _12598__674 (.L_HI(net674));
 sg13g2_tiehi _12597__675 (.L_HI(net675));
 sg13g2_tiehi _12596__676 (.L_HI(net676));
 sg13g2_tiehi _12595__677 (.L_HI(net677));
 sg13g2_tiehi _12594__678 (.L_HI(net678));
 sg13g2_tiehi _12593__679 (.L_HI(net679));
 sg13g2_tiehi _12592__680 (.L_HI(net680));
 sg13g2_tiehi _12591__681 (.L_HI(net681));
 sg13g2_tiehi _12590__682 (.L_HI(net682));
 sg13g2_tiehi _12589__683 (.L_HI(net683));
 sg13g2_tiehi _12917__684 (.L_HI(net684));
 sg13g2_tiehi _12588__685 (.L_HI(net685));
 sg13g2_tiehi _12586__686 (.L_HI(net686));
 sg13g2_tiehi _12585__687 (.L_HI(net687));
 sg13g2_tiehi _12584__688 (.L_HI(net688));
 sg13g2_tiehi _12583__689 (.L_HI(net689));
 sg13g2_tiehi _12582__690 (.L_HI(net690));
 sg13g2_tiehi _12581__691 (.L_HI(net691));
 sg13g2_tiehi _12580__692 (.L_HI(net692));
 sg13g2_tiehi _12579__693 (.L_HI(net693));
 sg13g2_tiehi _12578__694 (.L_HI(net694));
 sg13g2_tiehi _12577__695 (.L_HI(net695));
 sg13g2_tiehi _12576__696 (.L_HI(net696));
 sg13g2_tiehi _12575__697 (.L_HI(net697));
 sg13g2_tiehi _12574__698 (.L_HI(net698));
 sg13g2_tiehi _12573__699 (.L_HI(net699));
 sg13g2_tiehi _12572__700 (.L_HI(net700));
 sg13g2_tiehi _12571__701 (.L_HI(net701));
 sg13g2_tiehi _12916__702 (.L_HI(net702));
 sg13g2_tiehi _12915__703 (.L_HI(net703));
 sg13g2_tiehi _12914__704 (.L_HI(net704));
 sg13g2_tiehi _12913__705 (.L_HI(net705));
 sg13g2_tiehi _12912__706 (.L_HI(net706));
 sg13g2_tiehi _12911__707 (.L_HI(net707));
 sg13g2_tiehi _12910__708 (.L_HI(net708));
 sg13g2_tiehi _12909__709 (.L_HI(net709));
 sg13g2_tiehi _12908__710 (.L_HI(net710));
 sg13g2_tiehi _12907__711 (.L_HI(net711));
 sg13g2_tiehi _12906__712 (.L_HI(net712));
 sg13g2_tiehi _12905__713 (.L_HI(net713));
 sg13g2_tiehi _12904__714 (.L_HI(net714));
 sg13g2_tiehi _12903__715 (.L_HI(net715));
 sg13g2_tiehi _12902__716 (.L_HI(net716));
 sg13g2_tiehi _12901__717 (.L_HI(net717));
 sg13g2_tiehi _12900__718 (.L_HI(net718));
 sg13g2_tiehi _12899__719 (.L_HI(net719));
 sg13g2_tiehi _12898__720 (.L_HI(net720));
 sg13g2_tiehi _12897__721 (.L_HI(net721));
 sg13g2_tiehi _12896__722 (.L_HI(net722));
 sg13g2_tiehi _12895__723 (.L_HI(net723));
 sg13g2_tiehi _12894__724 (.L_HI(net724));
 sg13g2_tiehi _12893__725 (.L_HI(net725));
 sg13g2_tiehi _12892__726 (.L_HI(net726));
 sg13g2_tiehi _12747__727 (.L_HI(net727));
 sg13g2_tiehi _12943__728 (.L_HI(net728));
 sg13g2_tiehi _12945__729 (.L_HI(net729));
 sg13g2_tiehi _12946__730 (.L_HI(net730));
 sg13g2_tiehi _12947__731 (.L_HI(net731));
 sg13g2_tiehi _12948__732 (.L_HI(net732));
 sg13g2_tiehi _12949__733 (.L_HI(net733));
 sg13g2_tiehi _12950__734 (.L_HI(net734));
 sg13g2_tiehi _12951__735 (.L_HI(net735));
 sg13g2_tiehi _12952__736 (.L_HI(net736));
 sg13g2_tiehi _12953__737 (.L_HI(net737));
 sg13g2_tiehi _12954__738 (.L_HI(net738));
 sg13g2_tiehi _12955__739 (.L_HI(net739));
 sg13g2_tiehi _12956__740 (.L_HI(net740));
 sg13g2_tiehi _12957__741 (.L_HI(net741));
 sg13g2_tiehi _12958__742 (.L_HI(net742));
 sg13g2_tiehi _12959__743 (.L_HI(net743));
 sg13g2_tiehi _12960__744 (.L_HI(net744));
 sg13g2_tiehi _12961__745 (.L_HI(net745));
 sg13g2_tiehi _12962__746 (.L_HI(net746));
 sg13g2_tiehi _12963__747 (.L_HI(net747));
 sg13g2_tiehi _12964__748 (.L_HI(net748));
 sg13g2_tiehi _12965__749 (.L_HI(net749));
 sg13g2_tiehi _12966__750 (.L_HI(net750));
 sg13g2_tiehi _12967__751 (.L_HI(net751));
 sg13g2_tiehi _12968__752 (.L_HI(net752));
 sg13g2_tiehi _12969__753 (.L_HI(net753));
 sg13g2_tiehi _12970__754 (.L_HI(net754));
 sg13g2_tiehi _12971__755 (.L_HI(net755));
 sg13g2_tiehi _12972__756 (.L_HI(net756));
 sg13g2_tiehi _12973__757 (.L_HI(net757));
 sg13g2_tiehi _12974__758 (.L_HI(net758));
 sg13g2_tiehi _12891__759 (.L_HI(net759));
 sg13g2_tiehi _12890__760 (.L_HI(net760));
 sg13g2_tiehi _12548__761 (.L_HI(net761));
 sg13g2_tiehi _12547__762 (.L_HI(net762));
 sg13g2_tiehi _12546__763 (.L_HI(net763));
 sg13g2_tiehi _12545__764 (.L_HI(net764));
 sg13g2_tiehi _12544__765 (.L_HI(net765));
 sg13g2_tiehi _12543__766 (.L_HI(net766));
 sg13g2_tiehi _12542__767 (.L_HI(net767));
 sg13g2_tiehi _12541__768 (.L_HI(net768));
 sg13g2_tiehi _12540__769 (.L_HI(net769));
 sg13g2_tiehi _12539__770 (.L_HI(net770));
 sg13g2_tiehi _12538__771 (.L_HI(net771));
 sg13g2_tiehi _12537__772 (.L_HI(net772));
 sg13g2_tiehi _12536__773 (.L_HI(net773));
 sg13g2_tiehi _12535__774 (.L_HI(net774));
 sg13g2_tiehi _12534__775 (.L_HI(net775));
 sg13g2_tiehi _12533__776 (.L_HI(net776));
 sg13g2_tiehi _12532__777 (.L_HI(net777));
 sg13g2_tiehi _12531__778 (.L_HI(net778));
 sg13g2_tiehi _12530__779 (.L_HI(net779));
 sg13g2_tiehi _12529__780 (.L_HI(net780));
 sg13g2_tiehi _12528__781 (.L_HI(net781));
 sg13g2_tiehi _12527__782 (.L_HI(net782));
 sg13g2_tiehi _12526__783 (.L_HI(net783));
 sg13g2_tiehi _12525__784 (.L_HI(net784));
 sg13g2_tiehi _12524__785 (.L_HI(net785));
 sg13g2_tiehi _12523__786 (.L_HI(net786));
 sg13g2_tiehi _12522__787 (.L_HI(net787));
 sg13g2_tiehi _12975__788 (.L_HI(net788));
 sg13g2_tiehi _13007__789 (.L_HI(net789));
 sg13g2_tiehi _13008__790 (.L_HI(net790));
 sg13g2_tiehi _13009__791 (.L_HI(net791));
 sg13g2_tiehi _13010__792 (.L_HI(net792));
 sg13g2_tiehi _13011__793 (.L_HI(net793));
 sg13g2_tiehi _13012__794 (.L_HI(net794));
 sg13g2_tiehi _13013__795 (.L_HI(net795));
 sg13g2_tiehi _13014__796 (.L_HI(net796));
 sg13g2_tiehi _13015__797 (.L_HI(net797));
 sg13g2_tiehi _13016__798 (.L_HI(net798));
 sg13g2_tiehi _13017__799 (.L_HI(net799));
 sg13g2_tiehi _13018__800 (.L_HI(net800));
 sg13g2_tiehi _13019__801 (.L_HI(net801));
 sg13g2_tiehi _13020__802 (.L_HI(net802));
 sg13g2_tiehi _13021__803 (.L_HI(net803));
 sg13g2_tiehi _13022__804 (.L_HI(net804));
 sg13g2_tiehi _13023__805 (.L_HI(net805));
 sg13g2_tiehi _13024__806 (.L_HI(net806));
 sg13g2_tiehi _13025__807 (.L_HI(net807));
 sg13g2_tiehi _13026__808 (.L_HI(net808));
 sg13g2_tiehi _13027__809 (.L_HI(net809));
 sg13g2_tiehi _13028__810 (.L_HI(net810));
 sg13g2_tiehi _13029__811 (.L_HI(net811));
 sg13g2_tiehi _13030__812 (.L_HI(net812));
 sg13g2_tiehi _13031__813 (.L_HI(net813));
 sg13g2_tiehi _13032__814 (.L_HI(net814));
 sg13g2_tiehi _13033__815 (.L_HI(net815));
 sg13g2_tiehi _13034__816 (.L_HI(net816));
 sg13g2_tiehi _13035__817 (.L_HI(net817));
 sg13g2_tiehi _13036__818 (.L_HI(net818));
 sg13g2_tiehi _12521__819 (.L_HI(net819));
 sg13g2_tiehi _12520__820 (.L_HI(net820));
 sg13g2_tiehi _12519__821 (.L_HI(net821));
 sg13g2_tiehi _12518__822 (.L_HI(net822));
 sg13g2_tiehi _12517__823 (.L_HI(net823));
 sg13g2_tiehi _12516__824 (.L_HI(net824));
 sg13g2_tiehi _12515__825 (.L_HI(net825));
 sg13g2_tiehi _12514__826 (.L_HI(net826));
 sg13g2_tiehi _12513__827 (.L_HI(net827));
 sg13g2_tiehi _12512__828 (.L_HI(net828));
 sg13g2_tiehi _12511__829 (.L_HI(net829));
 sg13g2_tiehi _12510__830 (.L_HI(net830));
 sg13g2_tiehi _12509__831 (.L_HI(net831));
 sg13g2_tiehi _12508__832 (.L_HI(net832));
 sg13g2_tiehi _12507__833 (.L_HI(net833));
 sg13g2_tiehi _12506__834 (.L_HI(net834));
 sg13g2_tiehi _12505__835 (.L_HI(net835));
 sg13g2_tiehi _12504__836 (.L_HI(net836));
 sg13g2_tiehi _12503__837 (.L_HI(net837));
 sg13g2_tiehi _12502__838 (.L_HI(net838));
 sg13g2_tiehi _12501__839 (.L_HI(net839));
 sg13g2_tiehi _12500__840 (.L_HI(net840));
 sg13g2_tiehi _12499__841 (.L_HI(net841));
 sg13g2_tiehi _12498__842 (.L_HI(net842));
 sg13g2_tiehi _12497__843 (.L_HI(net843));
 sg13g2_tiehi _12496__844 (.L_HI(net844));
 sg13g2_tiehi _12495__845 (.L_HI(net845));
 sg13g2_tiehi _12494__846 (.L_HI(net846));
 sg13g2_tiehi _12493__847 (.L_HI(net847));
 sg13g2_tiehi _12492__848 (.L_HI(net848));
 sg13g2_tiehi _12491__849 (.L_HI(net849));
 sg13g2_tiehi _12490__850 (.L_HI(net850));
 sg13g2_tiehi _12489__851 (.L_HI(net851));
 sg13g2_tiehi _12488__852 (.L_HI(net852));
 sg13g2_tiehi _12487__853 (.L_HI(net853));
 sg13g2_tiehi _12486__854 (.L_HI(net854));
 sg13g2_tiehi _12485__855 (.L_HI(net855));
 sg13g2_tiehi _12484__856 (.L_HI(net856));
 sg13g2_tiehi _12483__857 (.L_HI(net857));
 sg13g2_tiehi _12482__858 (.L_HI(net858));
 sg13g2_tiehi _12481__859 (.L_HI(net859));
 sg13g2_tiehi _12480__860 (.L_HI(net860));
 sg13g2_tiehi _12479__861 (.L_HI(net861));
 sg13g2_tiehi _12478__862 (.L_HI(net862));
 sg13g2_tiehi _12477__863 (.L_HI(net863));
 sg13g2_tiehi _12476__864 (.L_HI(net864));
 sg13g2_tiehi _12475__865 (.L_HI(net865));
 sg13g2_tiehi _12474__866 (.L_HI(net866));
 sg13g2_tiehi _12473__867 (.L_HI(net867));
 sg13g2_tiehi _12472__868 (.L_HI(net868));
 sg13g2_tiehi _12471__869 (.L_HI(net869));
 sg13g2_tiehi _12470__870 (.L_HI(net870));
 sg13g2_tiehi _12469__871 (.L_HI(net871));
 sg13g2_tiehi _12468__872 (.L_HI(net872));
 sg13g2_tiehi _12467__873 (.L_HI(net873));
 sg13g2_tiehi _12466__874 (.L_HI(net874));
 sg13g2_tiehi _12465__875 (.L_HI(net875));
 sg13g2_tiehi _12464__876 (.L_HI(net876));
 sg13g2_tiehi _12463__877 (.L_HI(net877));
 sg13g2_tiehi _12462__878 (.L_HI(net878));
 sg13g2_tiehi _12461__879 (.L_HI(net879));
 sg13g2_tiehi _12460__880 (.L_HI(net880));
 sg13g2_tiehi _12459__881 (.L_HI(net881));
 sg13g2_tiehi _12458__882 (.L_HI(net882));
 sg13g2_tiehi _12457__883 (.L_HI(net883));
 sg13g2_tiehi _12456__884 (.L_HI(net884));
 sg13g2_tiehi _12455__885 (.L_HI(net885));
 sg13g2_tiehi _12454__886 (.L_HI(net886));
 sg13g2_tiehi _12453__887 (.L_HI(net887));
 sg13g2_tiehi _12452__888 (.L_HI(net888));
 sg13g2_tiehi _12451__889 (.L_HI(net889));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_1 _13983_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _13984_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _13985_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _13986_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _13987_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _13988_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _13989_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_2 _13990_ (.A(pwmpin),
    .X(uo_out[3]));
 sg13g2_buf_1 _13991_ (.A(net3049),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout2981 (.A(_04843_),
    .X(net2981));
 sg13g2_buf_2 fanout2982 (.A(_04843_),
    .X(net2982));
 sg13g2_buf_2 fanout2983 (.A(_04833_),
    .X(net2983));
 sg13g2_buf_2 fanout2984 (.A(_04833_),
    .X(net2984));
 sg13g2_buf_2 fanout2985 (.A(_04801_),
    .X(net2985));
 sg13g2_buf_2 fanout2986 (.A(_04801_),
    .X(net2986));
 sg13g2_buf_4 fanout2987 (.X(net2987),
    .A(_04790_));
 sg13g2_buf_2 fanout2988 (.A(_04790_),
    .X(net2988));
 sg13g2_buf_2 fanout2989 (.A(net2990),
    .X(net2989));
 sg13g2_buf_2 fanout2990 (.A(_04757_),
    .X(net2990));
 sg13g2_buf_2 fanout2991 (.A(net2992),
    .X(net2991));
 sg13g2_buf_4 fanout2992 (.X(net2992),
    .A(_04746_));
 sg13g2_buf_4 fanout2993 (.X(net2993),
    .A(_04734_));
 sg13g2_buf_2 fanout2994 (.A(_04734_),
    .X(net2994));
 sg13g2_buf_2 fanout2995 (.A(_04722_),
    .X(net2995));
 sg13g2_buf_2 fanout2996 (.A(_04722_),
    .X(net2996));
 sg13g2_buf_2 fanout2997 (.A(_04710_),
    .X(net2997));
 sg13g2_buf_2 fanout2998 (.A(_04710_),
    .X(net2998));
 sg13g2_buf_2 fanout2999 (.A(net3000),
    .X(net2999));
 sg13g2_buf_4 fanout3000 (.X(net3000),
    .A(_04698_));
 sg13g2_buf_4 fanout3001 (.X(net3001),
    .A(net3002));
 sg13g2_buf_4 fanout3002 (.X(net3002),
    .A(_04619_));
 sg13g2_buf_2 fanout3003 (.A(_04389_),
    .X(net3003));
 sg13g2_buf_2 fanout3004 (.A(_04389_),
    .X(net3004));
 sg13g2_buf_2 fanout3005 (.A(_04355_),
    .X(net3005));
 sg13g2_buf_2 fanout3006 (.A(_04355_),
    .X(net3006));
 sg13g2_buf_2 fanout3007 (.A(_04866_),
    .X(net3007));
 sg13g2_buf_4 fanout3008 (.X(net3008),
    .A(_04866_));
 sg13g2_buf_2 fanout3009 (.A(_04854_),
    .X(net3009));
 sg13g2_buf_2 fanout3010 (.A(_04854_),
    .X(net3010));
 sg13g2_buf_2 fanout3011 (.A(net3012),
    .X(net3011));
 sg13g2_buf_2 fanout3012 (.A(_04822_),
    .X(net3012));
 sg13g2_buf_2 fanout3013 (.A(net3014),
    .X(net3013));
 sg13g2_buf_4 fanout3014 (.X(net3014),
    .A(_04810_));
 sg13g2_buf_2 fanout3015 (.A(net3016),
    .X(net3015));
 sg13g2_buf_4 fanout3016 (.X(net3016),
    .A(_04780_));
 sg13g2_buf_2 fanout3017 (.A(_04768_),
    .X(net3017));
 sg13g2_buf_2 fanout3018 (.A(_04768_),
    .X(net3018));
 sg13g2_buf_4 fanout3019 (.X(net3019),
    .A(_04640_));
 sg13g2_buf_2 fanout3020 (.A(_04640_),
    .X(net3020));
 sg13g2_buf_2 fanout3021 (.A(_04597_),
    .X(net3021));
 sg13g2_buf_2 fanout3022 (.A(_04597_),
    .X(net3022));
 sg13g2_buf_2 fanout3023 (.A(_04572_),
    .X(net3023));
 sg13g2_buf_2 fanout3024 (.A(_04572_),
    .X(net3024));
 sg13g2_buf_2 fanout3025 (.A(net3026),
    .X(net3025));
 sg13g2_buf_2 fanout3026 (.A(_04543_),
    .X(net3026));
 sg13g2_buf_2 fanout3027 (.A(_04515_),
    .X(net3027));
 sg13g2_buf_2 fanout3028 (.A(_04515_),
    .X(net3028));
 sg13g2_buf_2 fanout3029 (.A(_04423_),
    .X(net3029));
 sg13g2_buf_2 fanout3030 (.A(_04423_),
    .X(net3030));
 sg13g2_buf_4 fanout3031 (.X(net3031),
    .A(_04686_));
 sg13g2_buf_2 fanout3032 (.A(_04686_),
    .X(net3032));
 sg13g2_buf_2 fanout3033 (.A(_04683_),
    .X(net3033));
 sg13g2_buf_2 fanout3034 (.A(_04683_),
    .X(net3034));
 sg13g2_buf_2 fanout3035 (.A(_04662_),
    .X(net3035));
 sg13g2_buf_2 fanout3036 (.A(_04662_),
    .X(net3036));
 sg13g2_buf_2 fanout3037 (.A(net3038),
    .X(net3037));
 sg13g2_buf_2 fanout3038 (.A(_04455_),
    .X(net3038));
 sg13g2_buf_2 fanout3039 (.A(net3040),
    .X(net3039));
 sg13g2_buf_2 fanout3040 (.A(_04326_),
    .X(net3040));
 sg13g2_buf_2 fanout3041 (.A(net3042),
    .X(net3041));
 sg13g2_buf_4 fanout3042 (.X(net3042),
    .A(_04298_));
 sg13g2_buf_4 fanout3043 (.X(net3043),
    .A(_04489_));
 sg13g2_buf_2 fanout3044 (.A(_04487_),
    .X(net3044));
 sg13g2_buf_2 fanout3045 (.A(_04487_),
    .X(net3045));
 sg13g2_buf_4 fanout3046 (.X(net3046),
    .A(_04263_));
 sg13g2_buf_2 fanout3047 (.A(_04263_),
    .X(net3047));
 sg13g2_buf_2 fanout3048 (.A(_03386_),
    .X(net3048));
 sg13g2_buf_2 fanout3049 (.A(net3049),
    .X(uio_oe[7]));
 sg13g2_buf_2 fanout3050 (.A(_02526_),
    .X(net3050));
 sg13g2_buf_2 fanout3051 (.A(_02526_),
    .X(net3051));
 sg13g2_buf_2 fanout3052 (.A(net3053),
    .X(net3052));
 sg13g2_buf_2 fanout3053 (.A(net3057),
    .X(net3053));
 sg13g2_buf_2 fanout3054 (.A(net3056),
    .X(net3054));
 sg13g2_buf_2 fanout3055 (.A(net3056),
    .X(net3055));
 sg13g2_buf_2 fanout3056 (.A(net3057),
    .X(net3056));
 sg13g2_buf_2 fanout3057 (.A(_05613_),
    .X(net3057));
 sg13g2_buf_2 fanout3058 (.A(net3059),
    .X(net3058));
 sg13g2_buf_4 fanout3059 (.X(net3059),
    .A(net3060));
 sg13g2_buf_4 fanout3060 (.X(net3060),
    .A(_05613_));
 sg13g2_buf_4 fanout3061 (.X(net3061),
    .A(_05006_));
 sg13g2_buf_2 fanout3062 (.A(net3063),
    .X(net3062));
 sg13g2_buf_2 fanout3063 (.A(_04960_),
    .X(net3063));
 sg13g2_buf_2 fanout3064 (.A(net3065),
    .X(net3064));
 sg13g2_buf_2 fanout3065 (.A(net3066),
    .X(net3065));
 sg13g2_buf_2 fanout3066 (.A(_04960_),
    .X(net3066));
 sg13g2_buf_2 fanout3067 (.A(net3069),
    .X(net3067));
 sg13g2_buf_4 fanout3068 (.X(net3068),
    .A(net3069));
 sg13g2_buf_2 fanout3069 (.A(_04960_),
    .X(net3069));
 sg13g2_buf_2 fanout3070 (.A(net3072),
    .X(net3070));
 sg13g2_buf_2 fanout3071 (.A(net3072),
    .X(net3071));
 sg13g2_buf_2 fanout3072 (.A(net3077),
    .X(net3072));
 sg13g2_buf_2 fanout3073 (.A(net3077),
    .X(net3073));
 sg13g2_buf_2 fanout3074 (.A(net3075),
    .X(net3074));
 sg13g2_buf_2 fanout3075 (.A(net3076),
    .X(net3075));
 sg13g2_buf_4 fanout3076 (.X(net3076),
    .A(net3077));
 sg13g2_buf_4 fanout3077 (.X(net3077),
    .A(_04929_));
 sg13g2_buf_2 fanout3078 (.A(net3082),
    .X(net3078));
 sg13g2_buf_2 fanout3079 (.A(net3081),
    .X(net3079));
 sg13g2_buf_2 fanout3080 (.A(net3081),
    .X(net3080));
 sg13g2_buf_2 fanout3081 (.A(net3082),
    .X(net3081));
 sg13g2_buf_2 fanout3082 (.A(_04869_),
    .X(net3082));
 sg13g2_buf_2 fanout3083 (.A(net3085),
    .X(net3083));
 sg13g2_buf_4 fanout3084 (.X(net3084),
    .A(net3085));
 sg13g2_buf_2 fanout3085 (.A(_04869_),
    .X(net3085));
 sg13g2_buf_2 fanout3086 (.A(net3089),
    .X(net3086));
 sg13g2_buf_2 fanout3087 (.A(net3088),
    .X(net3087));
 sg13g2_buf_2 fanout3088 (.A(net3089),
    .X(net3088));
 sg13g2_buf_2 fanout3089 (.A(_03436_),
    .X(net3089));
 sg13g2_buf_2 fanout3090 (.A(net3091),
    .X(net3090));
 sg13g2_buf_2 fanout3091 (.A(_03433_),
    .X(net3091));
 sg13g2_buf_2 fanout3092 (.A(net3097),
    .X(net3092));
 sg13g2_buf_2 fanout3093 (.A(net3097),
    .X(net3093));
 sg13g2_buf_2 fanout3094 (.A(net3097),
    .X(net3094));
 sg13g2_buf_1 fanout3095 (.A(net3096),
    .X(net3095));
 sg13g2_buf_4 fanout3096 (.X(net3096),
    .A(net3097));
 sg13g2_buf_2 fanout3097 (.A(_02569_),
    .X(net3097));
 sg13g2_buf_2 fanout3098 (.A(_02404_),
    .X(net3098));
 sg13g2_buf_2 fanout3099 (.A(_02404_),
    .X(net3099));
 sg13g2_buf_2 fanout3100 (.A(_05377_),
    .X(net3100));
 sg13g2_buf_1 fanout3101 (.A(_05377_),
    .X(net3101));
 sg13g2_buf_2 fanout3102 (.A(net3103),
    .X(net3102));
 sg13g2_buf_2 fanout3103 (.A(_05377_),
    .X(net3103));
 sg13g2_buf_2 fanout3104 (.A(net3106),
    .X(net3104));
 sg13g2_buf_1 fanout3105 (.A(net3106),
    .X(net3105));
 sg13g2_buf_4 fanout3106 (.X(net3106),
    .A(net3108));
 sg13g2_buf_4 fanout3107 (.X(net3107),
    .A(net3108));
 sg13g2_buf_2 fanout3108 (.A(_04067_),
    .X(net3108));
 sg13g2_buf_2 fanout3109 (.A(net3110),
    .X(net3109));
 sg13g2_buf_2 fanout3110 (.A(net3111),
    .X(net3110));
 sg13g2_buf_4 fanout3111 (.X(net3111),
    .A(net3113));
 sg13g2_buf_4 fanout3112 (.X(net3112),
    .A(net3113));
 sg13g2_buf_2 fanout3113 (.A(_04066_),
    .X(net3113));
 sg13g2_buf_2 fanout3114 (.A(net3116),
    .X(net3114));
 sg13g2_buf_4 fanout3115 (.X(net3115),
    .A(net3116));
 sg13g2_buf_2 fanout3116 (.A(_04062_),
    .X(net3116));
 sg13g2_buf_2 fanout3117 (.A(_02422_),
    .X(net3117));
 sg13g2_buf_2 fanout3118 (.A(net3119),
    .X(net3118));
 sg13g2_buf_2 fanout3119 (.A(_02413_),
    .X(net3119));
 sg13g2_buf_2 fanout3120 (.A(net3121),
    .X(net3120));
 sg13g2_buf_1 fanout3121 (.A(_02418_),
    .X(net3121));
 sg13g2_buf_2 fanout3122 (.A(_02412_),
    .X(net3122));
 sg13g2_buf_2 fanout3123 (.A(_02412_),
    .X(net3123));
 sg13g2_buf_4 fanout3124 (.X(net3124),
    .A(_03150_));
 sg13g2_buf_4 fanout3125 (.X(net3125),
    .A(_03149_));
 sg13g2_buf_2 fanout3126 (.A(net3128),
    .X(net3126));
 sg13g2_buf_1 fanout3127 (.A(net3128),
    .X(net3127));
 sg13g2_buf_2 fanout3128 (.A(_02417_),
    .X(net3128));
 sg13g2_buf_2 fanout3129 (.A(_04241_),
    .X(net3129));
 sg13g2_buf_2 fanout3130 (.A(net3131),
    .X(net3130));
 sg13g2_buf_2 fanout3131 (.A(net3132),
    .X(net3131));
 sg13g2_buf_2 fanout3132 (.A(net3133),
    .X(net3132));
 sg13g2_buf_2 fanout3133 (.A(_02516_),
    .X(net3133));
 sg13g2_buf_4 fanout3134 (.X(net3134),
    .A(_02505_));
 sg13g2_buf_2 fanout3135 (.A(net3136),
    .X(net3135));
 sg13g2_buf_2 fanout3136 (.A(net3139),
    .X(net3136));
 sg13g2_buf_2 fanout3137 (.A(net3138),
    .X(net3137));
 sg13g2_buf_1 fanout3138 (.A(net3139),
    .X(net3138));
 sg13g2_buf_4 fanout3139 (.X(net3139),
    .A(net3140));
 sg13g2_buf_4 fanout3140 (.X(net3140),
    .A(_02504_));
 sg13g2_buf_2 fanout3141 (.A(net3142),
    .X(net3141));
 sg13g2_buf_2 fanout3142 (.A(_02421_),
    .X(net3142));
 sg13g2_buf_8 fanout3143 (.A(net3148),
    .X(net3143));
 sg13g2_buf_4 fanout3144 (.X(net3144),
    .A(net3148));
 sg13g2_buf_8 fanout3145 (.A(net3148),
    .X(net3145));
 sg13g2_buf_4 fanout3146 (.X(net3146),
    .A(net3147));
 sg13g2_buf_4 fanout3147 (.X(net3147),
    .A(net3148));
 sg13g2_buf_8 fanout3148 (.A(_05560_),
    .X(net3148));
 sg13g2_buf_4 fanout3149 (.X(net3149),
    .A(net3150));
 sg13g2_buf_4 fanout3150 (.X(net3150),
    .A(net3154));
 sg13g2_buf_4 fanout3151 (.X(net3151),
    .A(net3154));
 sg13g2_buf_4 fanout3152 (.X(net3152),
    .A(net3153));
 sg13g2_buf_8 fanout3153 (.A(net3154),
    .X(net3153));
 sg13g2_buf_4 fanout3154 (.X(net3154),
    .A(_05039_));
 sg13g2_buf_8 fanout3155 (.A(net3157),
    .X(net3155));
 sg13g2_buf_2 fanout3156 (.A(net3157),
    .X(net3156));
 sg13g2_buf_4 fanout3157 (.X(net3157),
    .A(_05034_));
 sg13g2_buf_8 fanout3158 (.A(net3160),
    .X(net3158));
 sg13g2_buf_4 fanout3159 (.X(net3159),
    .A(net3160));
 sg13g2_buf_8 fanout3160 (.A(_05034_),
    .X(net3160));
 sg13g2_buf_8 fanout3161 (.A(net3162),
    .X(net3161));
 sg13g2_buf_8 fanout3162 (.A(net3166),
    .X(net3162));
 sg13g2_buf_4 fanout3163 (.X(net3163),
    .A(net3166));
 sg13g2_buf_4 fanout3164 (.X(net3164),
    .A(net3165));
 sg13g2_buf_8 fanout3165 (.A(net3166),
    .X(net3165));
 sg13g2_buf_4 fanout3166 (.X(net3166),
    .A(_05029_));
 sg13g2_buf_8 fanout3167 (.A(_04997_),
    .X(net3167));
 sg13g2_buf_4 fanout3168 (.X(net3168),
    .A(_04997_));
 sg13g2_buf_4 fanout3169 (.X(net3169),
    .A(net3172));
 sg13g2_buf_4 fanout3170 (.X(net3170),
    .A(net3171));
 sg13g2_buf_4 fanout3171 (.X(net3171),
    .A(net3172));
 sg13g2_buf_4 fanout3172 (.X(net3172),
    .A(_04997_));
 sg13g2_buf_8 fanout3173 (.A(net3178),
    .X(net3173));
 sg13g2_buf_2 fanout3174 (.A(net3178),
    .X(net3174));
 sg13g2_buf_8 fanout3175 (.A(net3178),
    .X(net3175));
 sg13g2_buf_4 fanout3176 (.X(net3176),
    .A(net3177));
 sg13g2_buf_4 fanout3177 (.X(net3177),
    .A(net3178));
 sg13g2_buf_8 fanout3178 (.A(_04992_),
    .X(net3178));
 sg13g2_buf_8 fanout3179 (.A(net3184),
    .X(net3179));
 sg13g2_buf_4 fanout3180 (.X(net3180),
    .A(net3184));
 sg13g2_buf_4 fanout3181 (.X(net3181),
    .A(net3184));
 sg13g2_buf_4 fanout3182 (.X(net3182),
    .A(net3183));
 sg13g2_buf_4 fanout3183 (.X(net3183),
    .A(net3184));
 sg13g2_buf_8 fanout3184 (.A(_04986_),
    .X(net3184));
 sg13g2_buf_4 fanout3185 (.X(net3185),
    .A(net3186));
 sg13g2_buf_8 fanout3186 (.A(net3190),
    .X(net3186));
 sg13g2_buf_4 fanout3187 (.X(net3187),
    .A(net3190));
 sg13g2_buf_4 fanout3188 (.X(net3188),
    .A(net3189));
 sg13g2_buf_8 fanout3189 (.A(net3190),
    .X(net3189));
 sg13g2_buf_4 fanout3190 (.X(net3190),
    .A(_04955_));
 sg13g2_buf_4 fanout3191 (.X(net3191),
    .A(net3192));
 sg13g2_buf_4 fanout3192 (.X(net3192),
    .A(net3193));
 sg13g2_buf_4 fanout3193 (.X(net3193),
    .A(_04924_));
 sg13g2_buf_8 fanout3194 (.A(net3196),
    .X(net3194));
 sg13g2_buf_4 fanout3195 (.X(net3195),
    .A(net3196));
 sg13g2_buf_8 fanout3196 (.A(_04924_),
    .X(net3196));
 sg13g2_buf_8 fanout3197 (.A(_04918_),
    .X(net3197));
 sg13g2_buf_4 fanout3198 (.X(net3198),
    .A(_04918_));
 sg13g2_buf_4 fanout3199 (.X(net3199),
    .A(net3202));
 sg13g2_buf_4 fanout3200 (.X(net3200),
    .A(net3201));
 sg13g2_buf_4 fanout3201 (.X(net3201),
    .A(net3202));
 sg13g2_buf_4 fanout3202 (.X(net3202),
    .A(_04918_));
 sg13g2_buf_8 fanout3203 (.A(net3208),
    .X(net3203));
 sg13g2_buf_4 fanout3204 (.X(net3204),
    .A(net3207));
 sg13g2_buf_4 fanout3205 (.X(net3205),
    .A(net3207));
 sg13g2_buf_4 fanout3206 (.X(net3206),
    .A(net3207));
 sg13g2_buf_4 fanout3207 (.X(net3207),
    .A(net3208));
 sg13g2_buf_4 fanout3208 (.X(net3208),
    .A(_04911_));
 sg13g2_buf_8 fanout3209 (.A(net3210),
    .X(net3209));
 sg13g2_buf_8 fanout3210 (.A(net3214),
    .X(net3210));
 sg13g2_buf_4 fanout3211 (.X(net3211),
    .A(net3214));
 sg13g2_buf_2 fanout3212 (.A(net3213),
    .X(net3212));
 sg13g2_buf_8 fanout3213 (.A(net3214),
    .X(net3213));
 sg13g2_buf_8 fanout3214 (.A(_04905_),
    .X(net3214));
 sg13g2_buf_4 fanout3215 (.X(net3215),
    .A(net3216));
 sg13g2_buf_8 fanout3216 (.A(_04898_),
    .X(net3216));
 sg13g2_buf_4 fanout3217 (.X(net3217),
    .A(net3218));
 sg13g2_buf_8 fanout3218 (.A(net3219),
    .X(net3218));
 sg13g2_buf_8 fanout3219 (.A(_04898_),
    .X(net3219));
 sg13g2_buf_8 fanout3220 (.A(net3225),
    .X(net3220));
 sg13g2_buf_4 fanout3221 (.X(net3221),
    .A(net3224));
 sg13g2_buf_4 fanout3222 (.X(net3222),
    .A(net3224));
 sg13g2_buf_4 fanout3223 (.X(net3223),
    .A(net3224));
 sg13g2_buf_8 fanout3224 (.A(net3225),
    .X(net3224));
 sg13g2_buf_4 fanout3225 (.X(net3225),
    .A(_04125_));
 sg13g2_buf_4 fanout3226 (.X(net3226),
    .A(net3227));
 sg13g2_buf_8 fanout3227 (.A(_05565_),
    .X(net3227));
 sg13g2_buf_4 fanout3228 (.X(net3228),
    .A(net3229));
 sg13g2_buf_8 fanout3229 (.A(net3230),
    .X(net3229));
 sg13g2_buf_8 fanout3230 (.A(_05565_),
    .X(net3230));
 sg13g2_buf_4 fanout3231 (.X(net3231),
    .A(net3233));
 sg13g2_buf_1 fanout3232 (.A(net3233),
    .X(net3232));
 sg13g2_buf_1 fanout3233 (.A(net3234),
    .X(net3233));
 sg13g2_buf_2 fanout3234 (.A(net3235),
    .X(net3234));
 sg13g2_buf_4 fanout3235 (.X(net3235),
    .A(net3236));
 sg13g2_buf_2 fanout3236 (.A(_02508_),
    .X(net3236));
 sg13g2_buf_4 fanout3237 (.X(net3237),
    .A(net3238));
 sg13g2_buf_4 fanout3238 (.X(net3238),
    .A(net3239));
 sg13g2_buf_2 fanout3239 (.A(_05572_),
    .X(net3239));
 sg13g2_buf_4 fanout3240 (.X(net3240),
    .A(_05572_));
 sg13g2_buf_2 fanout3241 (.A(net3242),
    .X(net3241));
 sg13g2_buf_2 fanout3242 (.A(net3243),
    .X(net3242));
 sg13g2_buf_2 fanout3243 (.A(_05571_),
    .X(net3243));
 sg13g2_buf_4 fanout3244 (.X(net3244),
    .A(_05571_));
 sg13g2_buf_4 fanout3245 (.X(net3245),
    .A(net3252));
 sg13g2_buf_2 fanout3246 (.A(net3252),
    .X(net3246));
 sg13g2_buf_4 fanout3247 (.X(net3247),
    .A(net3252));
 sg13g2_buf_4 fanout3248 (.X(net3248),
    .A(net3250));
 sg13g2_buf_4 fanout3249 (.X(net3249),
    .A(net3250));
 sg13g2_buf_2 fanout3250 (.A(net3251),
    .X(net3250));
 sg13g2_buf_2 fanout3251 (.A(net3252),
    .X(net3251));
 sg13g2_buf_2 fanout3252 (.A(_05059_),
    .X(net3252));
 sg13g2_buf_2 fanout3253 (.A(net3260),
    .X(net3253));
 sg13g2_buf_4 fanout3254 (.X(net3254),
    .A(net3260));
 sg13g2_buf_2 fanout3255 (.A(net3256),
    .X(net3255));
 sg13g2_buf_2 fanout3256 (.A(net3257),
    .X(net3256));
 sg13g2_buf_2 fanout3257 (.A(net3260),
    .X(net3257));
 sg13g2_buf_4 fanout3258 (.X(net3258),
    .A(net3259));
 sg13g2_buf_4 fanout3259 (.X(net3259),
    .A(net3260));
 sg13g2_buf_2 fanout3260 (.A(_05045_),
    .X(net3260));
 sg13g2_buf_2 fanout3261 (.A(net3264),
    .X(net3261));
 sg13g2_buf_2 fanout3262 (.A(net3264),
    .X(net3262));
 sg13g2_buf_1 fanout3263 (.A(net3264),
    .X(net3263));
 sg13g2_buf_1 fanout3264 (.A(net3265),
    .X(net3264));
 sg13g2_buf_2 fanout3265 (.A(net3267),
    .X(net3265));
 sg13g2_buf_2 fanout3266 (.A(net3267),
    .X(net3266));
 sg13g2_buf_2 fanout3267 (.A(_03747_),
    .X(net3267));
 sg13g2_buf_2 fanout3268 (.A(net3269),
    .X(net3268));
 sg13g2_buf_4 fanout3269 (.X(net3269),
    .A(_03746_));
 sg13g2_buf_2 fanout3270 (.A(net3272),
    .X(net3270));
 sg13g2_buf_1 fanout3271 (.A(net3272),
    .X(net3271));
 sg13g2_buf_2 fanout3272 (.A(net3273),
    .X(net3272));
 sg13g2_buf_2 fanout3273 (.A(_03691_),
    .X(net3273));
 sg13g2_buf_2 fanout3274 (.A(net3275),
    .X(net3274));
 sg13g2_buf_2 fanout3275 (.A(net3276),
    .X(net3275));
 sg13g2_buf_2 fanout3276 (.A(_03690_),
    .X(net3276));
 sg13g2_buf_2 fanout3277 (.A(_03690_),
    .X(net3277));
 sg13g2_buf_2 fanout3278 (.A(_03690_),
    .X(net3278));
 sg13g2_buf_2 fanout3279 (.A(net3283),
    .X(net3279));
 sg13g2_buf_1 fanout3280 (.A(net3283),
    .X(net3280));
 sg13g2_buf_2 fanout3281 (.A(net3282),
    .X(net3281));
 sg13g2_buf_2 fanout3282 (.A(net3283),
    .X(net3282));
 sg13g2_buf_2 fanout3283 (.A(net3284),
    .X(net3283));
 sg13g2_buf_2 fanout3284 (.A(_03680_),
    .X(net3284));
 sg13g2_buf_2 fanout3285 (.A(net3287),
    .X(net3285));
 sg13g2_buf_1 fanout3286 (.A(net3287),
    .X(net3286));
 sg13g2_buf_2 fanout3287 (.A(net3288),
    .X(net3287));
 sg13g2_buf_2 fanout3288 (.A(_03679_),
    .X(net3288));
 sg13g2_buf_4 fanout3289 (.X(net3289),
    .A(net3290));
 sg13g2_buf_2 fanout3290 (.A(_02500_),
    .X(net3290));
 sg13g2_buf_2 fanout3291 (.A(net3292),
    .X(net3291));
 sg13g2_buf_2 fanout3292 (.A(net3293),
    .X(net3292));
 sg13g2_buf_1 fanout3293 (.A(net3297),
    .X(net3293));
 sg13g2_buf_4 fanout3294 (.X(net3294),
    .A(net3297));
 sg13g2_buf_2 fanout3295 (.A(net3297),
    .X(net3295));
 sg13g2_buf_2 fanout3296 (.A(net3297),
    .X(net3296));
 sg13g2_buf_2 fanout3297 (.A(_02500_),
    .X(net3297));
 sg13g2_buf_2 fanout3298 (.A(net3301),
    .X(net3298));
 sg13g2_buf_2 fanout3299 (.A(net3300),
    .X(net3299));
 sg13g2_buf_2 fanout3300 (.A(net3301),
    .X(net3300));
 sg13g2_buf_2 fanout3301 (.A(net3302),
    .X(net3301));
 sg13g2_buf_2 fanout3302 (.A(net3307),
    .X(net3302));
 sg13g2_buf_2 fanout3303 (.A(net3304),
    .X(net3303));
 sg13g2_buf_2 fanout3304 (.A(net3307),
    .X(net3304));
 sg13g2_buf_2 fanout3305 (.A(net3307),
    .X(net3305));
 sg13g2_buf_1 fanout3306 (.A(net3307),
    .X(net3306));
 sg13g2_buf_1 fanout3307 (.A(_02475_),
    .X(net3307));
 sg13g2_buf_4 fanout3308 (.X(net3308),
    .A(net3309));
 sg13g2_buf_4 fanout3309 (.X(net3309),
    .A(_05046_));
 sg13g2_buf_4 fanout3310 (.X(net3310),
    .A(_04265_));
 sg13g2_buf_2 fanout3311 (.A(_04265_),
    .X(net3311));
 sg13g2_buf_2 fanout3312 (.A(net3313),
    .X(net3312));
 sg13g2_buf_2 fanout3313 (.A(_04264_),
    .X(net3313));
 sg13g2_buf_2 fanout3314 (.A(net3315),
    .X(net3314));
 sg13g2_buf_4 fanout3315 (.X(net3315),
    .A(net3316));
 sg13g2_buf_4 fanout3316 (.X(net3316),
    .A(net3318));
 sg13g2_buf_4 fanout3317 (.X(net3317),
    .A(net3318));
 sg13g2_buf_4 fanout3318 (.X(net3318),
    .A(_04121_));
 sg13g2_buf_4 fanout3319 (.X(net3319),
    .A(_04078_));
 sg13g2_buf_2 fanout3320 (.A(_04078_),
    .X(net3320));
 sg13g2_buf_8 fanout3321 (.A(net3325),
    .X(net3321));
 sg13g2_buf_8 fanout3322 (.A(net3325),
    .X(net3322));
 sg13g2_buf_4 fanout3323 (.X(net3323),
    .A(net3324));
 sg13g2_buf_2 fanout3324 (.A(net3325),
    .X(net3324));
 sg13g2_buf_4 fanout3325 (.X(net3325),
    .A(_04077_));
 sg13g2_buf_4 fanout3326 (.X(net3326),
    .A(_03101_));
 sg13g2_buf_4 fanout3327 (.X(net3327),
    .A(_03014_));
 sg13g2_buf_8 fanout3328 (.A(_02842_),
    .X(net3328));
 sg13g2_buf_8 fanout3329 (.A(_02759_),
    .X(net3329));
 sg13g2_buf_4 fanout3330 (.X(net3330),
    .A(_02663_));
 sg13g2_buf_4 fanout3331 (.X(net3331),
    .A(net3334));
 sg13g2_buf_4 fanout3332 (.X(net3332),
    .A(net3334));
 sg13g2_buf_4 fanout3333 (.X(net3333),
    .A(net3334));
 sg13g2_buf_4 fanout3334 (.X(net3334),
    .A(_02442_));
 sg13g2_buf_4 fanout3335 (.X(net3335),
    .A(_02441_));
 sg13g2_buf_2 fanout3336 (.A(_02441_),
    .X(net3336));
 sg13g2_buf_4 fanout3337 (.X(net3337),
    .A(_04285_));
 sg13g2_buf_2 fanout3338 (.A(_04285_),
    .X(net3338));
 sg13g2_buf_2 fanout3339 (.A(net3340),
    .X(net3339));
 sg13g2_buf_2 fanout3340 (.A(net3343),
    .X(net3340));
 sg13g2_buf_2 fanout3341 (.A(net3342),
    .X(net3341));
 sg13g2_buf_2 fanout3342 (.A(net3343),
    .X(net3342));
 sg13g2_buf_2 fanout3343 (.A(_04129_),
    .X(net3343));
 sg13g2_buf_2 fanout3344 (.A(net3346),
    .X(net3344));
 sg13g2_buf_2 fanout3345 (.A(net3346),
    .X(net3345));
 sg13g2_buf_2 fanout3346 (.A(net3347),
    .X(net3346));
 sg13g2_buf_2 fanout3347 (.A(_04129_),
    .X(net3347));
 sg13g2_buf_2 fanout3348 (.A(net3354),
    .X(net3348));
 sg13g2_buf_2 fanout3349 (.A(net3351),
    .X(net3349));
 sg13g2_buf_1 fanout3350 (.A(net3351),
    .X(net3350));
 sg13g2_buf_2 fanout3351 (.A(net3354),
    .X(net3351));
 sg13g2_buf_2 fanout3352 (.A(net3353),
    .X(net3352));
 sg13g2_buf_2 fanout3353 (.A(net3354),
    .X(net3353));
 sg13g2_buf_2 fanout3354 (.A(_04128_),
    .X(net3354));
 sg13g2_buf_2 fanout3355 (.A(net3356),
    .X(net3355));
 sg13g2_buf_4 fanout3356 (.X(net3356),
    .A(_04115_));
 sg13g2_buf_4 fanout3357 (.X(net3357),
    .A(net3358));
 sg13g2_buf_4 fanout3358 (.X(net3358),
    .A(_04114_));
 sg13g2_buf_2 fanout3359 (.A(net3360),
    .X(net3359));
 sg13g2_buf_2 fanout3360 (.A(_03668_),
    .X(net3360));
 sg13g2_buf_2 fanout3361 (.A(_03667_),
    .X(net3361));
 sg13g2_buf_2 fanout3362 (.A(net3363),
    .X(net3362));
 sg13g2_buf_2 fanout3363 (.A(net3364),
    .X(net3363));
 sg13g2_buf_2 fanout3364 (.A(net3365),
    .X(net3364));
 sg13g2_buf_4 fanout3365 (.X(net3365),
    .A(_03654_));
 sg13g2_buf_4 fanout3366 (.X(net3366),
    .A(net3367));
 sg13g2_buf_2 fanout3367 (.A(_02444_),
    .X(net3367));
 sg13g2_buf_4 fanout3368 (.X(net3368),
    .A(_02444_));
 sg13g2_buf_4 fanout3369 (.X(net3369),
    .A(net3370));
 sg13g2_buf_4 fanout3370 (.X(net3370),
    .A(_02443_));
 sg13g2_buf_2 fanout3371 (.A(net3373),
    .X(net3371));
 sg13g2_buf_1 fanout3372 (.A(net3373),
    .X(net3372));
 sg13g2_buf_4 fanout3373 (.X(net3373),
    .A(_04287_));
 sg13g2_buf_2 fanout3374 (.A(_04287_),
    .X(net3374));
 sg13g2_buf_2 fanout3375 (.A(_04287_),
    .X(net3375));
 sg13g2_buf_2 fanout3376 (.A(net3377),
    .X(net3376));
 sg13g2_buf_2 fanout3377 (.A(net3378),
    .X(net3377));
 sg13g2_buf_2 fanout3378 (.A(_04284_),
    .X(net3378));
 sg13g2_buf_2 fanout3379 (.A(net3382),
    .X(net3379));
 sg13g2_buf_1 fanout3380 (.A(net3382),
    .X(net3380));
 sg13g2_buf_2 fanout3381 (.A(net3382),
    .X(net3381));
 sg13g2_buf_2 fanout3382 (.A(_04065_),
    .X(net3382));
 sg13g2_buf_4 fanout3383 (.X(net3383),
    .A(_04065_));
 sg13g2_buf_1 fanout3384 (.A(_04065_),
    .X(net3384));
 sg13g2_buf_4 fanout3385 (.X(net3385),
    .A(_03659_));
 sg13g2_buf_8 fanout3386 (.A(_02482_),
    .X(net3386));
 sg13g2_buf_4 fanout3387 (.X(net3387),
    .A(net3389));
 sg13g2_buf_2 fanout3388 (.A(net3389),
    .X(net3388));
 sg13g2_buf_4 fanout3389 (.X(net3389),
    .A(_02472_));
 sg13g2_buf_2 fanout3390 (.A(net3391),
    .X(net3390));
 sg13g2_buf_2 fanout3391 (.A(_02431_),
    .X(net3391));
 sg13g2_buf_2 fanout3392 (.A(_02431_),
    .X(net3392));
 sg13g2_buf_4 fanout3393 (.X(net3393),
    .A(net3395));
 sg13g2_buf_4 fanout3394 (.X(net3394),
    .A(net3395));
 sg13g2_buf_2 fanout3395 (.A(_02431_),
    .X(net3395));
 sg13g2_buf_8 fanout3396 (.A(_01786_),
    .X(net3396));
 sg13g2_buf_2 fanout3397 (.A(_01786_),
    .X(net3397));
 sg13g2_buf_4 fanout3398 (.X(net3398),
    .A(net3400));
 sg13g2_buf_4 fanout3399 (.X(net3399),
    .A(net3400));
 sg13g2_buf_4 fanout3400 (.X(net3400),
    .A(_01786_));
 sg13g2_buf_2 fanout3401 (.A(net3402),
    .X(net3401));
 sg13g2_buf_2 fanout3402 (.A(net3403),
    .X(net3402));
 sg13g2_buf_2 fanout3403 (.A(net3404),
    .X(net3403));
 sg13g2_buf_2 fanout3404 (.A(net3405),
    .X(net3404));
 sg13g2_buf_4 fanout3405 (.X(net3405),
    .A(_01766_));
 sg13g2_buf_4 fanout3406 (.X(net3406),
    .A(net3407));
 sg13g2_buf_4 fanout3407 (.X(net3407),
    .A(_01765_));
 sg13g2_buf_4 fanout3408 (.X(net3408),
    .A(net3409));
 sg13g2_buf_4 fanout3409 (.X(net3409),
    .A(_04251_));
 sg13g2_buf_2 fanout3410 (.A(net3412),
    .X(net3410));
 sg13g2_buf_2 fanout3411 (.A(net3412),
    .X(net3411));
 sg13g2_buf_2 fanout3412 (.A(_04250_),
    .X(net3412));
 sg13g2_buf_2 fanout3413 (.A(net3415),
    .X(net3413));
 sg13g2_buf_4 fanout3414 (.X(net3414),
    .A(net3415));
 sg13g2_buf_2 fanout3415 (.A(_04064_),
    .X(net3415));
 sg13g2_buf_2 fanout3416 (.A(_02713_),
    .X(net3416));
 sg13g2_buf_2 fanout3417 (.A(_02539_),
    .X(net3417));
 sg13g2_buf_2 fanout3418 (.A(net3419),
    .X(net3418));
 sg13g2_buf_2 fanout3419 (.A(net3420),
    .X(net3419));
 sg13g2_buf_1 fanout3420 (.A(net3421),
    .X(net3420));
 sg13g2_buf_1 fanout3421 (.A(net3425),
    .X(net3421));
 sg13g2_buf_2 fanout3422 (.A(net3425),
    .X(net3422));
 sg13g2_buf_4 fanout3423 (.X(net3423),
    .A(net3425));
 sg13g2_buf_4 fanout3424 (.X(net3424),
    .A(net3425));
 sg13g2_buf_4 fanout3425 (.X(net3425),
    .A(_02471_));
 sg13g2_buf_8 fanout3426 (.A(net3429),
    .X(net3426));
 sg13g2_buf_4 fanout3427 (.X(net3427),
    .A(net3429));
 sg13g2_buf_4 fanout3428 (.X(net3428),
    .A(net3429));
 sg13g2_buf_8 fanout3429 (.A(_02462_),
    .X(net3429));
 sg13g2_buf_4 fanout3430 (.X(net3430),
    .A(_02459_));
 sg13g2_buf_2 fanout3431 (.A(_02459_),
    .X(net3431));
 sg13g2_buf_4 fanout3432 (.X(net3432),
    .A(net3434));
 sg13g2_buf_4 fanout3433 (.X(net3433),
    .A(net3434));
 sg13g2_buf_4 fanout3434 (.X(net3434),
    .A(_02459_));
 sg13g2_buf_2 fanout3435 (.A(net3437),
    .X(net3435));
 sg13g2_buf_2 fanout3436 (.A(net3438),
    .X(net3436));
 sg13g2_buf_1 fanout3437 (.A(net3438),
    .X(net3437));
 sg13g2_buf_4 fanout3438 (.X(net3438),
    .A(_02430_));
 sg13g2_buf_2 fanout3439 (.A(net3440),
    .X(net3439));
 sg13g2_buf_4 fanout3440 (.X(net3440),
    .A(_01783_));
 sg13g2_buf_8 fanout3441 (.A(_01782_),
    .X(net3441));
 sg13g2_buf_2 fanout3442 (.A(_01782_),
    .X(net3442));
 sg13g2_buf_4 fanout3443 (.X(net3443),
    .A(net3445));
 sg13g2_buf_4 fanout3444 (.X(net3444),
    .A(net3445));
 sg13g2_buf_4 fanout3445 (.X(net3445),
    .A(_01782_));
 sg13g2_buf_4 fanout3446 (.X(net3446),
    .A(net3447));
 sg13g2_buf_4 fanout3447 (.X(net3447),
    .A(_01780_));
 sg13g2_buf_2 fanout3448 (.A(_01763_),
    .X(net3448));
 sg13g2_buf_4 fanout3449 (.X(net3449),
    .A(_01763_));
 sg13g2_buf_2 fanout3450 (.A(net3451),
    .X(net3450));
 sg13g2_buf_4 fanout3451 (.X(net3451),
    .A(_01758_));
 sg13g2_buf_2 fanout3452 (.A(net3455),
    .X(net3452));
 sg13g2_buf_2 fanout3453 (.A(net3455),
    .X(net3453));
 sg13g2_buf_2 fanout3454 (.A(net3455),
    .X(net3454));
 sg13g2_buf_2 fanout3455 (.A(_04254_),
    .X(net3455));
 sg13g2_buf_2 fanout3456 (.A(net3457),
    .X(net3456));
 sg13g2_buf_4 fanout3457 (.X(net3457),
    .A(_02705_));
 sg13g2_buf_2 fanout3458 (.A(_02541_),
    .X(net3458));
 sg13g2_buf_2 fanout3459 (.A(_02509_),
    .X(net3459));
 sg13g2_buf_4 fanout3460 (.X(net3460),
    .A(net3461));
 sg13g2_buf_4 fanout3461 (.X(net3461),
    .A(net3463));
 sg13g2_buf_4 fanout3462 (.X(net3462),
    .A(net3463));
 sg13g2_buf_4 fanout3463 (.X(net3463),
    .A(_02453_));
 sg13g2_buf_4 fanout3464 (.X(net3464),
    .A(net3465));
 sg13g2_buf_4 fanout3465 (.X(net3465),
    .A(net3468));
 sg13g2_buf_4 fanout3466 (.X(net3466),
    .A(net3468));
 sg13g2_buf_4 fanout3467 (.X(net3467),
    .A(net3468));
 sg13g2_buf_8 fanout3468 (.A(_02450_),
    .X(net3468));
 sg13g2_buf_4 fanout3469 (.X(net3469),
    .A(net3470));
 sg13g2_buf_4 fanout3470 (.X(net3470),
    .A(net3473));
 sg13g2_buf_4 fanout3471 (.X(net3471),
    .A(net3472));
 sg13g2_buf_4 fanout3472 (.X(net3472),
    .A(net3473));
 sg13g2_buf_8 fanout3473 (.A(_02449_),
    .X(net3473));
 sg13g2_buf_4 fanout3474 (.X(net3474),
    .A(net3475));
 sg13g2_buf_2 fanout3475 (.A(net3476),
    .X(net3475));
 sg13g2_buf_2 fanout3476 (.A(net3483),
    .X(net3476));
 sg13g2_buf_4 fanout3477 (.X(net3477),
    .A(net3483));
 sg13g2_buf_4 fanout3478 (.X(net3478),
    .A(net3483));
 sg13g2_buf_2 fanout3479 (.A(net3483),
    .X(net3479));
 sg13g2_buf_4 fanout3480 (.X(net3480),
    .A(net3481));
 sg13g2_buf_4 fanout3481 (.X(net3481),
    .A(net3482));
 sg13g2_buf_4 fanout3482 (.X(net3482),
    .A(net3483));
 sg13g2_buf_4 fanout3483 (.X(net3483),
    .A(_02448_));
 sg13g2_buf_2 fanout3484 (.A(net3486),
    .X(net3484));
 sg13g2_buf_4 fanout3485 (.X(net3485),
    .A(net3486));
 sg13g2_buf_4 fanout3486 (.X(net3486),
    .A(net3510));
 sg13g2_buf_4 fanout3487 (.X(net3487),
    .A(net3489));
 sg13g2_buf_2 fanout3488 (.A(net3489),
    .X(net3488));
 sg13g2_buf_2 fanout3489 (.A(net3510),
    .X(net3489));
 sg13g2_buf_2 fanout3490 (.A(net3492),
    .X(net3490));
 sg13g2_buf_2 fanout3491 (.A(net3492),
    .X(net3491));
 sg13g2_buf_2 fanout3492 (.A(net3498),
    .X(net3492));
 sg13g2_buf_4 fanout3493 (.X(net3493),
    .A(net3498));
 sg13g2_buf_2 fanout3494 (.A(net3495),
    .X(net3494));
 sg13g2_buf_2 fanout3495 (.A(net3498),
    .X(net3495));
 sg13g2_buf_4 fanout3496 (.X(net3496),
    .A(net3497));
 sg13g2_buf_4 fanout3497 (.X(net3497),
    .A(net3498));
 sg13g2_buf_2 fanout3498 (.A(net3510),
    .X(net3498));
 sg13g2_buf_4 fanout3499 (.X(net3499),
    .A(net3500));
 sg13g2_buf_4 fanout3500 (.X(net3500),
    .A(net3504));
 sg13g2_buf_4 fanout3501 (.X(net3501),
    .A(net3504));
 sg13g2_buf_2 fanout3502 (.A(net3504),
    .X(net3502));
 sg13g2_buf_4 fanout3503 (.X(net3503),
    .A(net3504));
 sg13g2_buf_2 fanout3504 (.A(net3510),
    .X(net3504));
 sg13g2_buf_2 fanout3505 (.A(net3506),
    .X(net3505));
 sg13g2_buf_2 fanout3506 (.A(net3510),
    .X(net3506));
 sg13g2_buf_4 fanout3507 (.X(net3507),
    .A(net3509));
 sg13g2_buf_2 fanout3508 (.A(net3509),
    .X(net3508));
 sg13g2_buf_2 fanout3509 (.A(net3510),
    .X(net3509));
 sg13g2_buf_4 fanout3510 (.X(net3510),
    .A(_02448_));
 sg13g2_buf_8 fanout3511 (.A(net3516),
    .X(net3511));
 sg13g2_buf_4 fanout3512 (.X(net3512),
    .A(net3516));
 sg13g2_buf_4 fanout3513 (.X(net3513),
    .A(net3516));
 sg13g2_buf_4 fanout3514 (.X(net3514),
    .A(net3515));
 sg13g2_buf_4 fanout3515 (.X(net3515),
    .A(net3516));
 sg13g2_buf_8 fanout3516 (.A(_02447_),
    .X(net3516));
 sg13g2_buf_4 fanout3517 (.X(net3517),
    .A(net3520));
 sg13g2_buf_4 fanout3518 (.X(net3518),
    .A(net3520));
 sg13g2_buf_4 fanout3519 (.X(net3519),
    .A(net3520));
 sg13g2_buf_4 fanout3520 (.X(net3520),
    .A(_02446_));
 sg13g2_buf_4 fanout3521 (.X(net3521),
    .A(net3523));
 sg13g2_buf_4 fanout3522 (.X(net3522),
    .A(net3523));
 sg13g2_buf_4 fanout3523 (.X(net3523),
    .A(net3528));
 sg13g2_buf_4 fanout3524 (.X(net3524),
    .A(net3528));
 sg13g2_buf_2 fanout3525 (.A(net3528),
    .X(net3525));
 sg13g2_buf_2 fanout3526 (.A(net3527),
    .X(net3526));
 sg13g2_buf_4 fanout3527 (.X(net3527),
    .A(net3528));
 sg13g2_buf_2 fanout3528 (.A(_02446_),
    .X(net3528));
 sg13g2_buf_2 fanout3529 (.A(net3535),
    .X(net3529));
 sg13g2_buf_4 fanout3530 (.X(net3530),
    .A(net3535));
 sg13g2_buf_4 fanout3531 (.X(net3531),
    .A(net3534));
 sg13g2_buf_4 fanout3532 (.X(net3532),
    .A(net3533));
 sg13g2_buf_2 fanout3533 (.A(net3534),
    .X(net3533));
 sg13g2_buf_2 fanout3534 (.A(net3535),
    .X(net3534));
 sg13g2_buf_4 fanout3535 (.X(net3535),
    .A(_02445_));
 sg13g2_buf_2 fanout3536 (.A(net3539),
    .X(net3536));
 sg13g2_buf_1 fanout3537 (.A(net3539),
    .X(net3537));
 sg13g2_buf_4 fanout3538 (.X(net3538),
    .A(net3539));
 sg13g2_buf_2 fanout3539 (.A(net3553),
    .X(net3539));
 sg13g2_buf_2 fanout3540 (.A(net3541),
    .X(net3540));
 sg13g2_buf_4 fanout3541 (.X(net3541),
    .A(net3545));
 sg13g2_buf_2 fanout3542 (.A(net3543),
    .X(net3542));
 sg13g2_buf_2 fanout3543 (.A(net3544),
    .X(net3543));
 sg13g2_buf_4 fanout3544 (.X(net3544),
    .A(net3545));
 sg13g2_buf_2 fanout3545 (.A(net3553),
    .X(net3545));
 sg13g2_buf_4 fanout3546 (.X(net3546),
    .A(net3549));
 sg13g2_buf_4 fanout3547 (.X(net3547),
    .A(net3549));
 sg13g2_buf_2 fanout3548 (.A(net3549),
    .X(net3548));
 sg13g2_buf_2 fanout3549 (.A(net3553),
    .X(net3549));
 sg13g2_buf_2 fanout3550 (.A(net3552),
    .X(net3550));
 sg13g2_buf_4 fanout3551 (.X(net3551),
    .A(net3552));
 sg13g2_buf_2 fanout3552 (.A(net3553),
    .X(net3552));
 sg13g2_buf_4 fanout3553 (.X(net3553),
    .A(_02445_));
 sg13g2_buf_4 fanout3554 (.X(net3554),
    .A(net3568));
 sg13g2_buf_2 fanout3555 (.A(net3568),
    .X(net3555));
 sg13g2_buf_4 fanout3556 (.X(net3556),
    .A(net3558));
 sg13g2_buf_4 fanout3557 (.X(net3557),
    .A(net3558));
 sg13g2_buf_4 fanout3558 (.X(net3558),
    .A(net3568));
 sg13g2_buf_4 fanout3559 (.X(net3559),
    .A(net3560));
 sg13g2_buf_4 fanout3560 (.X(net3560),
    .A(net3567));
 sg13g2_buf_4 fanout3561 (.X(net3561),
    .A(net3563));
 sg13g2_buf_4 fanout3562 (.X(net3562),
    .A(net3567));
 sg13g2_buf_2 fanout3563 (.A(net3567),
    .X(net3563));
 sg13g2_buf_4 fanout3564 (.X(net3564),
    .A(net3566));
 sg13g2_buf_4 fanout3565 (.X(net3565),
    .A(net3566));
 sg13g2_buf_4 fanout3566 (.X(net3566),
    .A(net3567));
 sg13g2_buf_4 fanout3567 (.X(net3567),
    .A(net3568));
 sg13g2_buf_8 fanout3568 (.A(_01784_),
    .X(net3568));
 sg13g2_buf_4 fanout3569 (.X(net3569),
    .A(_01781_));
 sg13g2_buf_4 fanout3570 (.X(net3570),
    .A(net3571));
 sg13g2_buf_4 fanout3571 (.X(net3571),
    .A(net3572));
 sg13g2_buf_8 fanout3572 (.A(_01773_),
    .X(net3572));
 sg13g2_buf_4 fanout3573 (.X(net3573),
    .A(_01772_));
 sg13g2_buf_4 fanout3574 (.X(net3574),
    .A(net3584));
 sg13g2_buf_4 fanout3575 (.X(net3575),
    .A(net3576));
 sg13g2_buf_2 fanout3576 (.A(net3577),
    .X(net3576));
 sg13g2_buf_2 fanout3577 (.A(net3584),
    .X(net3577));
 sg13g2_buf_4 fanout3578 (.X(net3578),
    .A(net3579));
 sg13g2_buf_4 fanout3579 (.X(net3579),
    .A(net3584));
 sg13g2_buf_4 fanout3580 (.X(net3580),
    .A(net3582));
 sg13g2_buf_4 fanout3581 (.X(net3581),
    .A(net3582));
 sg13g2_buf_2 fanout3582 (.A(net3583),
    .X(net3582));
 sg13g2_buf_2 fanout3583 (.A(net3584),
    .X(net3583));
 sg13g2_buf_4 fanout3584 (.X(net3584),
    .A(_01769_));
 sg13g2_buf_4 fanout3585 (.X(net3585),
    .A(net3586));
 sg13g2_buf_4 fanout3586 (.X(net3586),
    .A(net3589));
 sg13g2_buf_4 fanout3587 (.X(net3587),
    .A(net3588));
 sg13g2_buf_2 fanout3588 (.A(net3589),
    .X(net3588));
 sg13g2_buf_4 fanout3589 (.X(net3589),
    .A(net3615));
 sg13g2_buf_4 fanout3590 (.X(net3590),
    .A(net3592));
 sg13g2_buf_2 fanout3591 (.A(net3592),
    .X(net3591));
 sg13g2_buf_4 fanout3592 (.X(net3592),
    .A(net3597));
 sg13g2_buf_4 fanout3593 (.X(net3593),
    .A(net3596));
 sg13g2_buf_4 fanout3594 (.X(net3594),
    .A(net3596));
 sg13g2_buf_2 fanout3595 (.A(net3596),
    .X(net3595));
 sg13g2_buf_4 fanout3596 (.X(net3596),
    .A(net3597));
 sg13g2_buf_2 fanout3597 (.A(net3615),
    .X(net3597));
 sg13g2_buf_2 fanout3598 (.A(net3606),
    .X(net3598));
 sg13g2_buf_2 fanout3599 (.A(net3606),
    .X(net3599));
 sg13g2_buf_4 fanout3600 (.X(net3600),
    .A(net3606));
 sg13g2_buf_2 fanout3601 (.A(net3605),
    .X(net3601));
 sg13g2_buf_2 fanout3602 (.A(net3605),
    .X(net3602));
 sg13g2_buf_4 fanout3603 (.X(net3603),
    .A(net3605));
 sg13g2_buf_2 fanout3604 (.A(net3605),
    .X(net3604));
 sg13g2_buf_2 fanout3605 (.A(net3606),
    .X(net3605));
 sg13g2_buf_2 fanout3606 (.A(net3615),
    .X(net3606));
 sg13g2_buf_2 fanout3607 (.A(net3608),
    .X(net3607));
 sg13g2_buf_4 fanout3608 (.X(net3608),
    .A(net3614));
 sg13g2_buf_2 fanout3609 (.A(net3611),
    .X(net3609));
 sg13g2_buf_1 fanout3610 (.A(net3611),
    .X(net3610));
 sg13g2_buf_2 fanout3611 (.A(net3613),
    .X(net3611));
 sg13g2_buf_2 fanout3612 (.A(net3613),
    .X(net3612));
 sg13g2_buf_2 fanout3613 (.A(net3614),
    .X(net3613));
 sg13g2_buf_2 fanout3614 (.A(net3615),
    .X(net3614));
 sg13g2_buf_4 fanout3615 (.X(net3615),
    .A(_01769_));
 sg13g2_buf_4 fanout3616 (.X(net3616),
    .A(net3618));
 sg13g2_buf_2 fanout3617 (.A(net3618),
    .X(net3617));
 sg13g2_buf_4 fanout3618 (.X(net3618),
    .A(net3619));
 sg13g2_buf_8 fanout3619 (.A(_01768_),
    .X(net3619));
 sg13g2_buf_4 fanout3620 (.X(net3620),
    .A(net3621));
 sg13g2_buf_4 fanout3621 (.X(net3621),
    .A(net3622));
 sg13g2_buf_4 fanout3622 (.X(net3622),
    .A(_01732_));
 sg13g2_buf_4 fanout3623 (.X(net3623),
    .A(_01730_));
 sg13g2_buf_4 fanout3624 (.X(net3624),
    .A(net3625));
 sg13g2_buf_4 fanout3625 (.X(net3625),
    .A(_01698_));
 sg13g2_buf_4 fanout3626 (.X(net3626),
    .A(net3627));
 sg13g2_buf_4 fanout3627 (.X(net3627),
    .A(_01691_));
 sg13g2_buf_4 fanout3628 (.X(net3628),
    .A(_01575_));
 sg13g2_buf_4 fanout3629 (.X(net3629),
    .A(net3630));
 sg13g2_buf_2 fanout3630 (.A(net3631),
    .X(net3630));
 sg13g2_buf_4 fanout3631 (.X(net3631),
    .A(net3634));
 sg13g2_buf_4 fanout3632 (.X(net3632),
    .A(net3633));
 sg13g2_buf_4 fanout3633 (.X(net3633),
    .A(net3634));
 sg13g2_buf_2 fanout3634 (.A(\cpu.mmode ),
    .X(net3634));
 sg13g2_buf_4 fanout3635 (.X(net3635),
    .A(net3637));
 sg13g2_buf_4 fanout3636 (.X(net3636),
    .A(net3637));
 sg13g2_buf_2 fanout3637 (.A(\cpu.mmode ),
    .X(net3637));
 sg13g2_buf_2 fanout3638 (.A(net3639),
    .X(net3638));
 sg13g2_buf_4 fanout3639 (.X(net3639),
    .A(_00059_));
 sg13g2_buf_2 fanout3640 (.A(_00059_),
    .X(net3640));
 sg13g2_buf_2 fanout3641 (.A(net3643),
    .X(net3641));
 sg13g2_buf_2 fanout3642 (.A(net3643),
    .X(net3642));
 sg13g2_buf_4 fanout3643 (.X(net3643),
    .A(net3644));
 sg13g2_buf_4 fanout3644 (.X(net3644),
    .A(\cpu.Bimm[12] ));
 sg13g2_buf_4 fanout3645 (.X(net3645),
    .A(net3646));
 sg13g2_buf_4 fanout3646 (.X(net3646),
    .A(net3653));
 sg13g2_buf_4 fanout3647 (.X(net3647),
    .A(net3653));
 sg13g2_buf_4 fanout3648 (.X(net3648),
    .A(net3652));
 sg13g2_buf_4 fanout3649 (.X(net3649),
    .A(net3651));
 sg13g2_buf_4 fanout3650 (.X(net3650),
    .A(net3651));
 sg13g2_buf_4 fanout3651 (.X(net3651),
    .A(net3652));
 sg13g2_buf_4 fanout3652 (.X(net3652),
    .A(net3653));
 sg13g2_buf_4 fanout3653 (.X(net3653),
    .A(\cpu.IR[20] ));
 sg13g2_buf_4 fanout3654 (.X(net3654),
    .A(net3655));
 sg13g2_buf_8 fanout3655 (.A(net3659),
    .X(net3655));
 sg13g2_buf_4 fanout3656 (.X(net3656),
    .A(net3658));
 sg13g2_buf_4 fanout3657 (.X(net3657),
    .A(net3659));
 sg13g2_buf_2 fanout3658 (.A(net3659),
    .X(net3658));
 sg13g2_buf_4 fanout3659 (.X(net3659),
    .A(\cpu.IR[17] ));
 sg13g2_buf_4 fanout3660 (.X(net3660),
    .A(net3661));
 sg13g2_buf_2 fanout3661 (.A(net3662),
    .X(net3661));
 sg13g2_buf_2 fanout3662 (.A(net3679),
    .X(net3662));
 sg13g2_buf_2 fanout3663 (.A(net3664),
    .X(net3663));
 sg13g2_buf_2 fanout3664 (.A(net3679),
    .X(net3664));
 sg13g2_buf_4 fanout3665 (.X(net3665),
    .A(net3679));
 sg13g2_buf_2 fanout3666 (.A(net3667),
    .X(net3666));
 sg13g2_buf_2 fanout3667 (.A(net3668),
    .X(net3667));
 sg13g2_buf_2 fanout3668 (.A(net3669),
    .X(net3668));
 sg13g2_buf_4 fanout3669 (.X(net3669),
    .A(net3679));
 sg13g2_buf_2 fanout3670 (.A(net3673),
    .X(net3670));
 sg13g2_buf_2 fanout3671 (.A(net3672),
    .X(net3671));
 sg13g2_buf_4 fanout3672 (.X(net3672),
    .A(net3673));
 sg13g2_buf_2 fanout3673 (.A(net3678),
    .X(net3673));
 sg13g2_buf_2 fanout3674 (.A(net3675),
    .X(net3674));
 sg13g2_buf_2 fanout3675 (.A(net3678),
    .X(net3675));
 sg13g2_buf_2 fanout3676 (.A(net3678),
    .X(net3676));
 sg13g2_buf_2 fanout3677 (.A(net3678),
    .X(net3677));
 sg13g2_buf_2 fanout3678 (.A(net3679),
    .X(net3678));
 sg13g2_buf_8 fanout3679 (.A(\cpu.IR[16] ),
    .X(net3679));
 sg13g2_buf_4 fanout3680 (.X(net3680),
    .A(net3685));
 sg13g2_buf_4 fanout3681 (.X(net3681),
    .A(net3684));
 sg13g2_buf_4 fanout3682 (.X(net3682),
    .A(net3683));
 sg13g2_buf_2 fanout3683 (.A(net3684),
    .X(net3683));
 sg13g2_buf_2 fanout3684 (.A(net3685),
    .X(net3684));
 sg13g2_buf_4 fanout3685 (.X(net3685),
    .A(\cpu.IR[15] ));
 sg13g2_buf_4 fanout3686 (.X(net3686),
    .A(net3687));
 sg13g2_buf_4 fanout3687 (.X(net3687),
    .A(net3688));
 sg13g2_buf_4 fanout3688 (.X(net3688),
    .A(\cpu.IR[15] ));
 sg13g2_buf_4 fanout3689 (.X(net3689),
    .A(net3690));
 sg13g2_buf_4 fanout3690 (.X(net3690),
    .A(net3693));
 sg13g2_buf_4 fanout3691 (.X(net3691),
    .A(net3693));
 sg13g2_buf_2 fanout3692 (.A(net3693),
    .X(net3692));
 sg13g2_buf_2 fanout3693 (.A(\cpu.IR[15] ),
    .X(net3693));
 sg13g2_buf_4 fanout3694 (.X(net3694),
    .A(\cpu.IR[14] ));
 sg13g2_buf_4 fanout3695 (.X(net3695),
    .A(net3697));
 sg13g2_buf_1 fanout3696 (.A(net3697),
    .X(net3696));
 sg13g2_buf_4 fanout3697 (.X(net3697),
    .A(\cpu.IR[13] ));
 sg13g2_buf_4 fanout3698 (.X(net3698),
    .A(\cpu.IR[13] ));
 sg13g2_buf_4 fanout3699 (.X(net3699),
    .A(\cpu.IR[12] ));
 sg13g2_buf_4 fanout3700 (.X(net3700),
    .A(net3703));
 sg13g2_buf_2 fanout3701 (.A(net3702),
    .X(net3701));
 sg13g2_buf_2 fanout3702 (.A(net3703),
    .X(net3702));
 sg13g2_buf_2 fanout3703 (.A(net3704),
    .X(net3703));
 sg13g2_buf_2 fanout3704 (.A(\cpu.opvalid ),
    .X(net3704));
 sg13g2_buf_4 fanout3705 (.X(net3705),
    .A(net3722));
 sg13g2_buf_2 fanout3706 (.A(net3722),
    .X(net3706));
 sg13g2_buf_4 fanout3707 (.X(net3707),
    .A(net3710));
 sg13g2_buf_4 fanout3708 (.X(net3708),
    .A(net3710));
 sg13g2_buf_4 fanout3709 (.X(net3709),
    .A(net3710));
 sg13g2_buf_2 fanout3710 (.A(net3712),
    .X(net3710));
 sg13g2_buf_4 fanout3711 (.X(net3711),
    .A(net3712));
 sg13g2_buf_2 fanout3712 (.A(net3722),
    .X(net3712));
 sg13g2_buf_4 fanout3713 (.X(net3713),
    .A(net3714));
 sg13g2_buf_4 fanout3714 (.X(net3714),
    .A(net3717));
 sg13g2_buf_4 fanout3715 (.X(net3715),
    .A(net3716));
 sg13g2_buf_4 fanout3716 (.X(net3716),
    .A(net3717));
 sg13g2_buf_4 fanout3717 (.X(net3717),
    .A(net3719));
 sg13g2_buf_4 fanout3718 (.X(net3718),
    .A(net3719));
 sg13g2_buf_4 fanout3719 (.X(net3719),
    .A(net3722));
 sg13g2_buf_4 fanout3720 (.X(net3720),
    .A(net3721));
 sg13g2_buf_4 fanout3721 (.X(net3721),
    .A(net3722));
 sg13g2_buf_8 fanout3722 (.A(_00027_),
    .X(net3722));
 sg13g2_buf_2 fanout3723 (.A(net3724),
    .X(net3723));
 sg13g2_buf_4 fanout3724 (.X(net3724),
    .A(_02707_));
 sg13g2_buf_2 fanout3725 (.A(net3726),
    .X(net3725));
 sg13g2_buf_1 fanout3726 (.A(net3727),
    .X(net3726));
 sg13g2_buf_4 fanout3727 (.X(net3727),
    .A(_02686_));
 sg13g2_buf_2 fanout3728 (.A(_02630_),
    .X(net3728));
 sg13g2_buf_4 fanout3729 (.X(net3729),
    .A(net3733));
 sg13g2_buf_1 fanout3730 (.A(net3733),
    .X(net3730));
 sg13g2_buf_2 fanout3731 (.A(net3733),
    .X(net3731));
 sg13g2_buf_1 fanout3732 (.A(net3733),
    .X(net3732));
 sg13g2_buf_1 fanout3733 (.A(_02588_),
    .X(net3733));
 sg13g2_buf_4 fanout3734 (.X(net3734),
    .A(net3737));
 sg13g2_buf_2 fanout3735 (.A(net3737),
    .X(net3735));
 sg13g2_buf_2 fanout3736 (.A(net3737),
    .X(net3736));
 sg13g2_buf_2 fanout3737 (.A(_02567_),
    .X(net3737));
 sg13g2_buf_4 fanout3738 (.X(net3738),
    .A(\uart0.urxsh[0] ));
 sg13g2_buf_2 fanout3739 (.A(\uart0.urxsh[0] ),
    .X(net3739));
 sg13g2_buf_2 fanout3740 (.A(net3742),
    .X(net3740));
 sg13g2_buf_1 fanout3741 (.A(net3742),
    .X(net3741));
 sg13g2_buf_2 fanout3742 (.A(net3749),
    .X(net3742));
 sg13g2_buf_2 fanout3743 (.A(net3748),
    .X(net3743));
 sg13g2_buf_2 fanout3744 (.A(net3748),
    .X(net3744));
 sg13g2_buf_2 fanout3745 (.A(net3747),
    .X(net3745));
 sg13g2_buf_2 fanout3746 (.A(net3747),
    .X(net3746));
 sg13g2_buf_2 fanout3747 (.A(net3748),
    .X(net3747));
 sg13g2_buf_2 fanout3748 (.A(net3749),
    .X(net3748));
 sg13g2_buf_2 fanout3749 (.A(net3798),
    .X(net3749));
 sg13g2_buf_2 fanout3750 (.A(net3752),
    .X(net3750));
 sg13g2_buf_2 fanout3751 (.A(net3752),
    .X(net3751));
 sg13g2_buf_2 fanout3752 (.A(net3760),
    .X(net3752));
 sg13g2_buf_2 fanout3753 (.A(net3755),
    .X(net3753));
 sg13g2_buf_2 fanout3754 (.A(net3755),
    .X(net3754));
 sg13g2_buf_2 fanout3755 (.A(net3760),
    .X(net3755));
 sg13g2_buf_2 fanout3756 (.A(net3757),
    .X(net3756));
 sg13g2_buf_2 fanout3757 (.A(net3759),
    .X(net3757));
 sg13g2_buf_1 fanout3758 (.A(net3759),
    .X(net3758));
 sg13g2_buf_4 fanout3759 (.X(net3759),
    .A(net3760));
 sg13g2_buf_2 fanout3760 (.A(net3798),
    .X(net3760));
 sg13g2_buf_2 fanout3761 (.A(net3763),
    .X(net3761));
 sg13g2_buf_4 fanout3762 (.X(net3762),
    .A(net3766));
 sg13g2_buf_2 fanout3763 (.A(net3766),
    .X(net3763));
 sg13g2_buf_2 fanout3764 (.A(net3766),
    .X(net3764));
 sg13g2_buf_2 fanout3765 (.A(net3766),
    .X(net3765));
 sg13g2_buf_1 fanout3766 (.A(net3778),
    .X(net3766));
 sg13g2_buf_4 fanout3767 (.X(net3767),
    .A(net3769));
 sg13g2_buf_4 fanout3768 (.X(net3768),
    .A(net3769));
 sg13g2_buf_1 fanout3769 (.A(net3771),
    .X(net3769));
 sg13g2_buf_4 fanout3770 (.X(net3770),
    .A(net3771));
 sg13g2_buf_2 fanout3771 (.A(net3778),
    .X(net3771));
 sg13g2_buf_2 fanout3772 (.A(net3776),
    .X(net3772));
 sg13g2_buf_1 fanout3773 (.A(net3776),
    .X(net3773));
 sg13g2_buf_4 fanout3774 (.X(net3774),
    .A(net3776));
 sg13g2_buf_1 fanout3775 (.A(net3776),
    .X(net3775));
 sg13g2_buf_1 fanout3776 (.A(net3778),
    .X(net3776));
 sg13g2_buf_4 fanout3777 (.X(net3777),
    .A(net3778));
 sg13g2_buf_2 fanout3778 (.A(net3798),
    .X(net3778));
 sg13g2_buf_2 fanout3779 (.A(net3780),
    .X(net3779));
 sg13g2_buf_2 fanout3780 (.A(net3798),
    .X(net3780));
 sg13g2_buf_2 fanout3781 (.A(net3786),
    .X(net3781));
 sg13g2_buf_2 fanout3782 (.A(net3786),
    .X(net3782));
 sg13g2_buf_2 fanout3783 (.A(net3785),
    .X(net3783));
 sg13g2_buf_2 fanout3784 (.A(net3785),
    .X(net3784));
 sg13g2_buf_4 fanout3785 (.X(net3785),
    .A(net3786));
 sg13g2_buf_1 fanout3786 (.A(net3797),
    .X(net3786));
 sg13g2_buf_2 fanout3787 (.A(net3788),
    .X(net3787));
 sg13g2_buf_1 fanout3788 (.A(net3797),
    .X(net3788));
 sg13g2_buf_2 fanout3789 (.A(net3791),
    .X(net3789));
 sg13g2_buf_1 fanout3790 (.A(net3791),
    .X(net3790));
 sg13g2_buf_2 fanout3791 (.A(net3797),
    .X(net3791));
 sg13g2_buf_2 fanout3792 (.A(net3793),
    .X(net3792));
 sg13g2_buf_2 fanout3793 (.A(net3796),
    .X(net3793));
 sg13g2_buf_2 fanout3794 (.A(net3795),
    .X(net3794));
 sg13g2_buf_2 fanout3795 (.A(net3796),
    .X(net3795));
 sg13g2_buf_2 fanout3796 (.A(net3797),
    .X(net3796));
 sg13g2_buf_2 fanout3797 (.A(net3798),
    .X(net3797));
 sg13g2_buf_4 fanout3798 (.X(net3798),
    .A(cclk));
 sg13g2_buf_4 fanout3799 (.X(net3799),
    .A(net3801));
 sg13g2_buf_2 fanout3800 (.A(net3801),
    .X(net3800));
 sg13g2_buf_2 fanout3801 (.A(net3802),
    .X(net3801));
 sg13g2_buf_2 fanout3802 (.A(net3812),
    .X(net3802));
 sg13g2_buf_2 fanout3803 (.A(net3805),
    .X(net3803));
 sg13g2_buf_2 fanout3804 (.A(net3808),
    .X(net3804));
 sg13g2_buf_1 fanout3805 (.A(net3808),
    .X(net3805));
 sg13g2_buf_2 fanout3806 (.A(net3807),
    .X(net3806));
 sg13g2_buf_4 fanout3807 (.X(net3807),
    .A(net3808));
 sg13g2_buf_2 fanout3808 (.A(net3812),
    .X(net3808));
 sg13g2_buf_2 fanout3809 (.A(net3811),
    .X(net3809));
 sg13g2_buf_2 fanout3810 (.A(net3811),
    .X(net3810));
 sg13g2_buf_2 fanout3811 (.A(net3812),
    .X(net3811));
 sg13g2_buf_2 fanout3812 (.A(net3870),
    .X(net3812));
 sg13g2_buf_2 fanout3813 (.A(net3815),
    .X(net3813));
 sg13g2_buf_2 fanout3814 (.A(net3815),
    .X(net3814));
 sg13g2_buf_2 fanout3815 (.A(net3823),
    .X(net3815));
 sg13g2_buf_2 fanout3816 (.A(net3823),
    .X(net3816));
 sg13g2_buf_2 fanout3817 (.A(net3823),
    .X(net3817));
 sg13g2_buf_2 fanout3818 (.A(net3819),
    .X(net3818));
 sg13g2_buf_2 fanout3819 (.A(net3822),
    .X(net3819));
 sg13g2_buf_2 fanout3820 (.A(net3821),
    .X(net3820));
 sg13g2_buf_2 fanout3821 (.A(net3822),
    .X(net3821));
 sg13g2_buf_2 fanout3822 (.A(net3823),
    .X(net3822));
 sg13g2_buf_2 fanout3823 (.A(net3870),
    .X(net3823));
 sg13g2_buf_2 fanout3824 (.A(net3833),
    .X(net3824));
 sg13g2_buf_2 fanout3825 (.A(net3833),
    .X(net3825));
 sg13g2_buf_2 fanout3826 (.A(net3827),
    .X(net3826));
 sg13g2_buf_2 fanout3827 (.A(net3833),
    .X(net3827));
 sg13g2_buf_2 fanout3828 (.A(net3829),
    .X(net3828));
 sg13g2_buf_2 fanout3829 (.A(net3832),
    .X(net3829));
 sg13g2_buf_2 fanout3830 (.A(net3832),
    .X(net3830));
 sg13g2_buf_2 fanout3831 (.A(net3832),
    .X(net3831));
 sg13g2_buf_4 fanout3832 (.X(net3832),
    .A(net3833));
 sg13g2_buf_1 fanout3833 (.A(net3870),
    .X(net3833));
 sg13g2_buf_2 fanout3834 (.A(net3838),
    .X(net3834));
 sg13g2_buf_1 fanout3835 (.A(net3838),
    .X(net3835));
 sg13g2_buf_2 fanout3836 (.A(net3837),
    .X(net3836));
 sg13g2_buf_2 fanout3837 (.A(net3838),
    .X(net3837));
 sg13g2_buf_2 fanout3838 (.A(net3839),
    .X(net3838));
 sg13g2_buf_2 fanout3839 (.A(net3870),
    .X(net3839));
 sg13g2_buf_2 fanout3840 (.A(net3850),
    .X(net3840));
 sg13g2_buf_2 fanout3841 (.A(net3850),
    .X(net3841));
 sg13g2_buf_2 fanout3842 (.A(net3844),
    .X(net3842));
 sg13g2_buf_2 fanout3843 (.A(net3844),
    .X(net3843));
 sg13g2_buf_2 fanout3844 (.A(net3850),
    .X(net3844));
 sg13g2_buf_2 fanout3845 (.A(net3846),
    .X(net3845));
 sg13g2_buf_2 fanout3846 (.A(net3849),
    .X(net3846));
 sg13g2_buf_2 fanout3847 (.A(net3849),
    .X(net3847));
 sg13g2_buf_2 fanout3848 (.A(net3849),
    .X(net3848));
 sg13g2_buf_2 fanout3849 (.A(net3850),
    .X(net3849));
 sg13g2_buf_2 fanout3850 (.A(net3870),
    .X(net3850));
 sg13g2_buf_2 fanout3851 (.A(net3855),
    .X(net3851));
 sg13g2_buf_2 fanout3852 (.A(net3855),
    .X(net3852));
 sg13g2_buf_2 fanout3853 (.A(net3855),
    .X(net3853));
 sg13g2_buf_2 fanout3854 (.A(net3855),
    .X(net3854));
 sg13g2_buf_2 fanout3855 (.A(net3869),
    .X(net3855));
 sg13g2_buf_2 fanout3856 (.A(net3857),
    .X(net3856));
 sg13g2_buf_2 fanout3857 (.A(net3860),
    .X(net3857));
 sg13g2_buf_2 fanout3858 (.A(net3860),
    .X(net3858));
 sg13g2_buf_2 fanout3859 (.A(net3860),
    .X(net3859));
 sg13g2_buf_2 fanout3860 (.A(net3869),
    .X(net3860));
 sg13g2_buf_2 fanout3861 (.A(net3862),
    .X(net3861));
 sg13g2_buf_2 fanout3862 (.A(net3866),
    .X(net3862));
 sg13g2_buf_2 fanout3863 (.A(net3865),
    .X(net3863));
 sg13g2_buf_2 fanout3864 (.A(net3865),
    .X(net3864));
 sg13g2_buf_2 fanout3865 (.A(net3866),
    .X(net3865));
 sg13g2_buf_2 fanout3866 (.A(net3869),
    .X(net3866));
 sg13g2_buf_2 fanout3867 (.A(net3868),
    .X(net3867));
 sg13g2_buf_2 fanout3868 (.A(net3869),
    .X(net3868));
 sg13g2_buf_2 fanout3869 (.A(net3870),
    .X(net3869));
 sg13g2_buf_8 fanout3870 (.A(cclk),
    .X(net3870));
 sg13g2_buf_2 fanout3871 (.A(net3872),
    .X(net3871));
 sg13g2_buf_4 fanout3872 (.X(net3872),
    .A(net3874));
 sg13g2_buf_2 fanout3873 (.A(net3874),
    .X(net3873));
 sg13g2_buf_2 fanout3874 (.A(net3876),
    .X(net3874));
 sg13g2_buf_2 fanout3875 (.A(net3876),
    .X(net3875));
 sg13g2_buf_4 fanout3876 (.X(net3876),
    .A(_03355_));
 sg13g2_buf_4 fanout3877 (.X(net3877),
    .A(net3880));
 sg13g2_buf_2 fanout3878 (.A(net3880),
    .X(net3878));
 sg13g2_buf_4 fanout3879 (.X(net3879),
    .A(net3880));
 sg13g2_buf_2 fanout3880 (.A(net3886),
    .X(net3880));
 sg13g2_buf_2 fanout3881 (.A(net3886),
    .X(net3881));
 sg13g2_buf_4 fanout3882 (.X(net3882),
    .A(net3883));
 sg13g2_buf_2 fanout3883 (.A(net3884),
    .X(net3883));
 sg13g2_buf_2 fanout3884 (.A(net3885),
    .X(net3884));
 sg13g2_buf_4 fanout3885 (.X(net3885),
    .A(net3886));
 sg13g2_buf_4 fanout3886 (.X(net3886),
    .A(_02591_));
 sg13g2_buf_2 fanout3887 (.A(net3890),
    .X(net3887));
 sg13g2_buf_2 fanout3888 (.A(net3890),
    .X(net3888));
 sg13g2_buf_2 fanout3889 (.A(net3890),
    .X(net3889));
 sg13g2_buf_2 fanout3890 (.A(net3891),
    .X(net3890));
 sg13g2_buf_2 fanout3891 (.A(net3898),
    .X(net3891));
 sg13g2_buf_2 fanout3892 (.A(net3893),
    .X(net3892));
 sg13g2_buf_2 fanout3893 (.A(net3898),
    .X(net3893));
 sg13g2_buf_2 fanout3894 (.A(net3896),
    .X(net3894));
 sg13g2_buf_2 fanout3895 (.A(net3896),
    .X(net3895));
 sg13g2_buf_2 fanout3896 (.A(net3897),
    .X(net3896));
 sg13g2_buf_2 fanout3897 (.A(net3898),
    .X(net3897));
 sg13g2_buf_4 fanout3898 (.X(net3898),
    .A(_02587_));
 sg13g2_buf_2 fanout3899 (.A(net3903),
    .X(net3899));
 sg13g2_buf_2 fanout3900 (.A(net3903),
    .X(net3900));
 sg13g2_buf_4 fanout3901 (.X(net3901),
    .A(net3902));
 sg13g2_buf_2 fanout3902 (.A(net3903),
    .X(net3902));
 sg13g2_buf_2 fanout3903 (.A(_02566_),
    .X(net3903));
 sg13g2_buf_4 fanout3904 (.X(net3904),
    .A(net3907));
 sg13g2_buf_1 fanout3905 (.A(net3907),
    .X(net3905));
 sg13g2_buf_2 fanout3906 (.A(net3907),
    .X(net3906));
 sg13g2_buf_2 fanout3907 (.A(_02552_),
    .X(net3907));
 sg13g2_buf_2 fanout3908 (.A(net3910),
    .X(net3908));
 sg13g2_buf_4 fanout3909 (.X(net3909),
    .A(net3910));
 sg13g2_buf_2 fanout3910 (.A(_02552_),
    .X(net3910));
 sg13g2_buf_2 fanout3911 (.A(net3913),
    .X(net3911));
 sg13g2_buf_1 fanout3912 (.A(net3913),
    .X(net3912));
 sg13g2_buf_2 fanout3913 (.A(net3914),
    .X(net3913));
 sg13g2_buf_2 fanout3914 (.A(net3920),
    .X(net3914));
 sg13g2_buf_2 fanout3915 (.A(net3917),
    .X(net3915));
 sg13g2_buf_2 fanout3916 (.A(net3917),
    .X(net3916));
 sg13g2_buf_2 fanout3917 (.A(net3920),
    .X(net3917));
 sg13g2_buf_2 fanout3918 (.A(net3920),
    .X(net3918));
 sg13g2_buf_2 fanout3919 (.A(net3920),
    .X(net3919));
 sg13g2_buf_2 fanout3920 (.A(_00545_),
    .X(net3920));
 sg13g2_buf_2 fanout3921 (.A(net3922),
    .X(net3921));
 sg13g2_buf_2 fanout3922 (.A(net3924),
    .X(net3922));
 sg13g2_buf_4 fanout3923 (.X(net3923),
    .A(net3924));
 sg13g2_buf_2 fanout3924 (.A(_00545_),
    .X(net3924));
 sg13g2_buf_2 fanout3925 (.A(\ckd[0] ),
    .X(net3925));
 sg13g2_buf_2 fanout3926 (.A(\jtag0.tapst[2] ),
    .X(net3926));
 sg13g2_buf_4 fanout3927 (.X(net3927),
    .A(\jtag0.tapst[0] ));
 sg13g2_buf_2 fanout3928 (.A(\jtag0.tapst[0] ),
    .X(net3928));
 sg13g2_buf_2 fanout3929 (.A(net3931),
    .X(net3929));
 sg13g2_buf_4 fanout3930 (.X(net3930),
    .A(net3931));
 sg13g2_buf_2 fanout3931 (.A(exintest),
    .X(net3931));
 sg13g2_buf_2 fanout3932 (.A(net3934),
    .X(net3932));
 sg13g2_buf_4 fanout3933 (.X(net3933),
    .A(net3934));
 sg13g2_buf_2 fanout3934 (.A(exintest),
    .X(net3934));
 sg13g2_buf_2 fanout3935 (.A(net3937),
    .X(net3935));
 sg13g2_buf_2 fanout3936 (.A(net3937),
    .X(net3936));
 sg13g2_buf_2 fanout3937 (.A(net3939),
    .X(net3937));
 sg13g2_buf_2 fanout3938 (.A(net3939),
    .X(net3938));
 sg13g2_buf_2 fanout3939 (.A(ui_in[0]),
    .X(net3939));
 sg13g2_buf_2 fanout3940 (.A(net3942),
    .X(net3940));
 sg13g2_buf_2 fanout3941 (.A(net3942),
    .X(net3941));
 sg13g2_buf_2 fanout3942 (.A(net3945),
    .X(net3942));
 sg13g2_buf_2 fanout3943 (.A(net3944),
    .X(net3943));
 sg13g2_buf_2 fanout3944 (.A(net3945),
    .X(net3944));
 sg13g2_buf_1 fanout3945 (.A(net3952),
    .X(net3945));
 sg13g2_buf_2 fanout3946 (.A(net3948),
    .X(net3946));
 sg13g2_buf_2 fanout3947 (.A(net3952),
    .X(net3947));
 sg13g2_buf_1 fanout3948 (.A(net3952),
    .X(net3948));
 sg13g2_buf_2 fanout3949 (.A(net3951),
    .X(net3949));
 sg13g2_buf_2 fanout3950 (.A(net3951),
    .X(net3950));
 sg13g2_buf_2 fanout3951 (.A(net3952),
    .X(net3951));
 sg13g2_buf_4 fanout3952 (.X(net3952),
    .A(ui_in[0]));
 sg13g2_buf_4 fanout3953 (.X(net3953),
    .A(net1));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _12450__17 (.L_HI(net17));
 sg13g2_buf_2 clkbuf_regs_1_clk (.A(jclk),
    .X(jclk_regs));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_0_jclk (.A(jclk),
    .X(clknet_0_jclk));
 sg13g2_buf_2 clkbuf_1_0__f_jclk (.A(clknet_0_jclk),
    .X(clknet_1_0__leaf_jclk));
 sg13g2_buf_2 clkbuf_1_1__f_jclk (.A(clknet_0_jclk),
    .X(clknet_1_1__leaf_jclk));
 sg13g2_buf_1 clkload1 (.A(clknet_1_1__leaf_jclk));
 sg13g2_buf_2 clkbuf_0_jclk_regs (.A(jclk_regs),
    .X(clknet_0_jclk_regs));
 sg13g2_buf_2 clkbuf_2_0__f_jclk_regs (.A(clknet_0_jclk_regs),
    .X(clknet_2_0__leaf_jclk_regs));
 sg13g2_buf_2 clkbuf_2_1__f_jclk_regs (.A(clknet_0_jclk_regs),
    .X(clknet_2_1__leaf_jclk_regs));
 sg13g2_buf_2 clkbuf_2_2__f_jclk_regs (.A(clknet_0_jclk_regs),
    .X(clknet_2_2__leaf_jclk_regs));
 sg13g2_buf_2 clkbuf_2_3__f_jclk_regs (.A(clknet_0_jclk_regs),
    .X(clknet_2_3__leaf_jclk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_jclk_regs));
 sg13g2_buf_2 clkbuf_0__02583_ (.A(_02583_),
    .X(clknet_0__02583_));
 sg13g2_buf_2 clkbuf_1_0__f__02583_ (.A(clknet_0__02583_),
    .X(clknet_1_0__leaf__02583_));
 sg13g2_buf_2 clkbuf_1_1__f__02583_ (.A(clknet_0__02583_),
    .X(clknet_1_1__leaf__02583_));
 sg13g2_buf_1 clkload3 (.A(clknet_1_0__leaf__02583_));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(delaynet_2_clk));
 sg13g2_buf_2 delaybuf_2_clk (.A(delaynet_2_clk),
    .X(clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00544_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold2 (.A(\xdi[13] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold3 (.A(_01151_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold4 (.A(\xdi[21] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold5 (.A(_01445_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold6 (.A(\xdi[7] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold7 (.A(_01145_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold8 (.A(\xdi[5] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold9 (.A(_01143_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold10 (.A(\xdi[4] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold11 (.A(\xdi[0] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold12 (.A(\xdi[2] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold13 (.A(_01140_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold14 (.A(\xdi[6] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold15 (.A(\xdi[3] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold16 (.A(\xdi[19] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold17 (.A(\xdi[10] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold18 (.A(_01148_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold19 (.A(\xdi[12] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold20 (.A(\xdi[11] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold21 (.A(\xdi[17] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold22 (.A(_01441_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold23 (.A(\xdi[23] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold24 (.A(_01447_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold25 (.A(\xdi[1] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold26 (.A(_01139_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold27 (.A(\xdi[9] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold28 (.A(_01147_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold29 (.A(\xdi[20] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold30 (.A(\xdi[15] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold31 (.A(_01153_),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold32 (.A(\xdi[16] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold33 (.A(\xdi[8] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold34 (.A(\xdi[18] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold35 (.A(_01442_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold36 (.A(\xdi[22] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold37 (.A(\xdi[14] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ckd[2] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold39 (.A(_00002_),
    .X(net928));
 sg13g2_antennanp ANTENNA_1 (.A(_02796_));
 sg13g2_antennanp ANTENNA_2 (.A(_02796_));
 sg13g2_antennanp ANTENNA_3 (.A(_02796_));
 sg13g2_antennanp ANTENNA_4 (.A(_02879_));
 sg13g2_antennanp ANTENNA_5 (.A(_02879_));
 sg13g2_antennanp ANTENNA_6 (.A(_02879_));
 sg13g2_antennanp ANTENNA_7 (.A(_02879_));
 sg13g2_antennanp ANTENNA_8 (.A(_02879_));
 sg13g2_antennanp ANTENNA_9 (.A(_03265_));
 sg13g2_antennanp ANTENNA_10 (.A(_03265_));
 sg13g2_antennanp ANTENNA_11 (.A(_03265_));
 sg13g2_antennanp ANTENNA_12 (.A(_03265_));
 sg13g2_antennanp ANTENNA_13 (.A(_04757_));
 sg13g2_antennanp ANTENNA_14 (.A(_04768_));
 sg13g2_antennanp ANTENNA_15 (.A(_04768_));
 sg13g2_antennanp ANTENNA_16 (.A(_04768_));
 sg13g2_antennanp ANTENNA_17 (.A(_04822_));
 sg13g2_antennanp ANTENNA_18 (.A(_04757_));
 sg13g2_antennanp ANTENNA_19 (.A(_04822_));
 sg13g2_antennanp ANTENNA_20 (.A(_04757_));
 sg13g2_antennanp ANTENNA_21 (.A(_04822_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_151 ();
 sg13g2_decap_4 FILLER_0_183 ();
 sg13g2_fill_1 FILLER_0_187 ();
 sg13g2_decap_4 FILLER_0_192 ();
 sg13g2_fill_1 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_decap_4 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_4 FILLER_0_234 ();
 sg13g2_fill_2 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_247 ();
 sg13g2_decap_4 FILLER_0_252 ();
 sg13g2_decap_4 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_4 FILLER_0_298 ();
 sg13g2_fill_1 FILLER_0_302 ();
 sg13g2_fill_2 FILLER_0_312 ();
 sg13g2_fill_1 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_fill_2 FILLER_0_417 ();
 sg13g2_fill_1 FILLER_0_419 ();
 sg13g2_decap_8 FILLER_0_432 ();
 sg13g2_decap_4 FILLER_0_439 ();
 sg13g2_decap_4 FILLER_0_469 ();
 sg13g2_fill_2 FILLER_0_473 ();
 sg13g2_decap_8 FILLER_0_501 ();
 sg13g2_decap_4 FILLER_0_508 ();
 sg13g2_fill_2 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_4 FILLER_0_547 ();
 sg13g2_fill_1 FILLER_0_551 ();
 sg13g2_fill_2 FILLER_0_562 ();
 sg13g2_fill_1 FILLER_0_564 ();
 sg13g2_decap_8 FILLER_0_579 ();
 sg13g2_decap_4 FILLER_0_586 ();
 sg13g2_fill_1 FILLER_0_590 ();
 sg13g2_decap_4 FILLER_0_601 ();
 sg13g2_fill_2 FILLER_0_605 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_fill_2 FILLER_0_680 ();
 sg13g2_fill_1 FILLER_0_682 ();
 sg13g2_fill_2 FILLER_0_693 ();
 sg13g2_fill_1 FILLER_0_695 ();
 sg13g2_fill_2 FILLER_0_723 ();
 sg13g2_fill_1 FILLER_0_725 ();
 sg13g2_decap_4 FILLER_0_752 ();
 sg13g2_fill_2 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_762 ();
 sg13g2_decap_4 FILLER_0_769 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_fill_1 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_4 FILLER_0_819 ();
 sg13g2_fill_1 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_fill_2 FILLER_0_835 ();
 sg13g2_fill_2 FILLER_0_847 ();
 sg13g2_fill_1 FILLER_0_849 ();
 sg13g2_decap_4 FILLER_0_854 ();
 sg13g2_fill_2 FILLER_0_858 ();
 sg13g2_decap_4 FILLER_0_873 ();
 sg13g2_fill_2 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_883 ();
 sg13g2_decap_8 FILLER_0_890 ();
 sg13g2_fill_1 FILLER_0_897 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_fill_2 FILLER_0_926 ();
 sg13g2_fill_1 FILLER_0_928 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_fill_2 FILLER_0_946 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_fill_1 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_970 ();
 sg13g2_decap_8 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_984 ();
 sg13g2_decap_8 FILLER_0_991 ();
 sg13g2_decap_8 FILLER_0_998 ();
 sg13g2_decap_8 FILLER_0_1005 ();
 sg13g2_decap_8 FILLER_0_1012 ();
 sg13g2_decap_8 FILLER_0_1019 ();
 sg13g2_decap_8 FILLER_0_1026 ();
 sg13g2_decap_8 FILLER_0_1033 ();
 sg13g2_decap_8 FILLER_0_1040 ();
 sg13g2_decap_8 FILLER_0_1047 ();
 sg13g2_decap_8 FILLER_0_1054 ();
 sg13g2_decap_8 FILLER_0_1061 ();
 sg13g2_decap_8 FILLER_0_1068 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_decap_8 FILLER_0_1103 ();
 sg13g2_decap_8 FILLER_0_1110 ();
 sg13g2_decap_8 FILLER_0_1117 ();
 sg13g2_decap_8 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1138 ();
 sg13g2_decap_8 FILLER_0_1145 ();
 sg13g2_decap_8 FILLER_0_1152 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1173 ();
 sg13g2_decap_8 FILLER_0_1180 ();
 sg13g2_decap_8 FILLER_0_1187 ();
 sg13g2_decap_8 FILLER_0_1194 ();
 sg13g2_decap_8 FILLER_0_1201 ();
 sg13g2_decap_8 FILLER_0_1208 ();
 sg13g2_decap_8 FILLER_0_1215 ();
 sg13g2_decap_8 FILLER_0_1222 ();
 sg13g2_decap_8 FILLER_0_1229 ();
 sg13g2_decap_8 FILLER_0_1236 ();
 sg13g2_decap_8 FILLER_0_1243 ();
 sg13g2_decap_8 FILLER_0_1250 ();
 sg13g2_decap_8 FILLER_0_1257 ();
 sg13g2_decap_8 FILLER_0_1264 ();
 sg13g2_decap_8 FILLER_0_1271 ();
 sg13g2_decap_8 FILLER_0_1278 ();
 sg13g2_decap_8 FILLER_0_1285 ();
 sg13g2_decap_8 FILLER_0_1292 ();
 sg13g2_decap_8 FILLER_0_1299 ();
 sg13g2_decap_8 FILLER_0_1306 ();
 sg13g2_fill_2 FILLER_0_1313 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_fill_2 FILLER_1_133 ();
 sg13g2_fill_1 FILLER_1_135 ();
 sg13g2_decap_4 FILLER_1_228 ();
 sg13g2_fill_1 FILLER_1_232 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_fill_2 FILLER_1_386 ();
 sg13g2_fill_1 FILLER_1_388 ();
 sg13g2_fill_2 FILLER_1_445 ();
 sg13g2_decap_4 FILLER_1_477 ();
 sg13g2_fill_1 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_decap_4 FILLER_1_647 ();
 sg13g2_fill_2 FILLER_1_655 ();
 sg13g2_fill_1 FILLER_1_657 ();
 sg13g2_fill_1 FILLER_1_668 ();
 sg13g2_decap_4 FILLER_1_731 ();
 sg13g2_decap_4 FILLER_1_743 ();
 sg13g2_fill_2 FILLER_1_793 ();
 sg13g2_fill_1 FILLER_1_795 ();
 sg13g2_fill_2 FILLER_1_866 ();
 sg13g2_fill_1 FILLER_1_930 ();
 sg13g2_fill_1 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_988 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1002 ();
 sg13g2_decap_8 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1016 ();
 sg13g2_decap_8 FILLER_1_1023 ();
 sg13g2_decap_8 FILLER_1_1030 ();
 sg13g2_decap_8 FILLER_1_1037 ();
 sg13g2_decap_8 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1051 ();
 sg13g2_decap_8 FILLER_1_1058 ();
 sg13g2_decap_8 FILLER_1_1065 ();
 sg13g2_decap_8 FILLER_1_1072 ();
 sg13g2_decap_8 FILLER_1_1079 ();
 sg13g2_decap_8 FILLER_1_1086 ();
 sg13g2_decap_8 FILLER_1_1093 ();
 sg13g2_decap_8 FILLER_1_1100 ();
 sg13g2_decap_8 FILLER_1_1107 ();
 sg13g2_decap_8 FILLER_1_1114 ();
 sg13g2_decap_8 FILLER_1_1121 ();
 sg13g2_decap_8 FILLER_1_1128 ();
 sg13g2_decap_8 FILLER_1_1135 ();
 sg13g2_decap_8 FILLER_1_1142 ();
 sg13g2_decap_8 FILLER_1_1149 ();
 sg13g2_decap_8 FILLER_1_1156 ();
 sg13g2_decap_8 FILLER_1_1163 ();
 sg13g2_decap_8 FILLER_1_1170 ();
 sg13g2_decap_8 FILLER_1_1177 ();
 sg13g2_decap_8 FILLER_1_1184 ();
 sg13g2_decap_8 FILLER_1_1191 ();
 sg13g2_decap_8 FILLER_1_1198 ();
 sg13g2_decap_8 FILLER_1_1205 ();
 sg13g2_decap_8 FILLER_1_1212 ();
 sg13g2_decap_8 FILLER_1_1219 ();
 sg13g2_decap_8 FILLER_1_1226 ();
 sg13g2_decap_8 FILLER_1_1233 ();
 sg13g2_decap_8 FILLER_1_1240 ();
 sg13g2_decap_8 FILLER_1_1247 ();
 sg13g2_decap_8 FILLER_1_1254 ();
 sg13g2_decap_8 FILLER_1_1261 ();
 sg13g2_decap_8 FILLER_1_1268 ();
 sg13g2_decap_8 FILLER_1_1275 ();
 sg13g2_decap_8 FILLER_1_1282 ();
 sg13g2_decap_8 FILLER_1_1289 ();
 sg13g2_decap_8 FILLER_1_1296 ();
 sg13g2_decap_8 FILLER_1_1303 ();
 sg13g2_decap_4 FILLER_1_1310 ();
 sg13g2_fill_1 FILLER_1_1314 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_4 FILLER_2_140 ();
 sg13g2_fill_2 FILLER_2_144 ();
 sg13g2_decap_4 FILLER_2_150 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_4 FILLER_2_224 ();
 sg13g2_fill_1 FILLER_2_228 ();
 sg13g2_fill_2 FILLER_2_276 ();
 sg13g2_fill_2 FILLER_2_287 ();
 sg13g2_fill_1 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_4 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_4 FILLER_2_366 ();
 sg13g2_decap_4 FILLER_2_396 ();
 sg13g2_fill_2 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_2 FILLER_2_420 ();
 sg13g2_fill_1 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_435 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_fill_1 FILLER_2_466 ();
 sg13g2_decap_4 FILLER_2_478 ();
 sg13g2_fill_2 FILLER_2_482 ();
 sg13g2_fill_2 FILLER_2_492 ();
 sg13g2_fill_1 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_499 ();
 sg13g2_decap_8 FILLER_2_506 ();
 sg13g2_decap_8 FILLER_2_513 ();
 sg13g2_decap_8 FILLER_2_520 ();
 sg13g2_decap_8 FILLER_2_527 ();
 sg13g2_decap_4 FILLER_2_534 ();
 sg13g2_fill_1 FILLER_2_542 ();
 sg13g2_decap_4 FILLER_2_553 ();
 sg13g2_fill_1 FILLER_2_557 ();
 sg13g2_fill_1 FILLER_2_584 ();
 sg13g2_decap_4 FILLER_2_599 ();
 sg13g2_fill_1 FILLER_2_603 ();
 sg13g2_fill_2 FILLER_2_614 ();
 sg13g2_fill_1 FILLER_2_616 ();
 sg13g2_fill_1 FILLER_2_621 ();
 sg13g2_decap_8 FILLER_2_626 ();
 sg13g2_decap_4 FILLER_2_633 ();
 sg13g2_decap_4 FILLER_2_673 ();
 sg13g2_fill_2 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_4 FILLER_2_710 ();
 sg13g2_decap_4 FILLER_2_750 ();
 sg13g2_fill_1 FILLER_2_758 ();
 sg13g2_decap_4 FILLER_2_779 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_4 FILLER_2_852 ();
 sg13g2_fill_1 FILLER_2_856 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_4 FILLER_2_914 ();
 sg13g2_fill_2 FILLER_2_918 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_4 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_965 ();
 sg13g2_decap_8 FILLER_2_972 ();
 sg13g2_decap_4 FILLER_2_979 ();
 sg13g2_decap_4 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_decap_8 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1036 ();
 sg13g2_decap_8 FILLER_2_1043 ();
 sg13g2_decap_8 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1057 ();
 sg13g2_decap_8 FILLER_2_1064 ();
 sg13g2_decap_8 FILLER_2_1071 ();
 sg13g2_decap_8 FILLER_2_1078 ();
 sg13g2_decap_8 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1092 ();
 sg13g2_decap_8 FILLER_2_1099 ();
 sg13g2_decap_8 FILLER_2_1106 ();
 sg13g2_decap_8 FILLER_2_1113 ();
 sg13g2_decap_8 FILLER_2_1120 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_8 FILLER_2_1134 ();
 sg13g2_decap_8 FILLER_2_1141 ();
 sg13g2_decap_8 FILLER_2_1148 ();
 sg13g2_decap_8 FILLER_2_1155 ();
 sg13g2_decap_8 FILLER_2_1162 ();
 sg13g2_decap_8 FILLER_2_1169 ();
 sg13g2_decap_8 FILLER_2_1176 ();
 sg13g2_decap_8 FILLER_2_1183 ();
 sg13g2_decap_8 FILLER_2_1190 ();
 sg13g2_decap_8 FILLER_2_1197 ();
 sg13g2_decap_8 FILLER_2_1204 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_decap_8 FILLER_2_1218 ();
 sg13g2_decap_8 FILLER_2_1225 ();
 sg13g2_decap_8 FILLER_2_1232 ();
 sg13g2_decap_8 FILLER_2_1239 ();
 sg13g2_decap_8 FILLER_2_1246 ();
 sg13g2_decap_8 FILLER_2_1253 ();
 sg13g2_decap_8 FILLER_2_1260 ();
 sg13g2_decap_8 FILLER_2_1267 ();
 sg13g2_decap_8 FILLER_2_1274 ();
 sg13g2_decap_8 FILLER_2_1281 ();
 sg13g2_decap_8 FILLER_2_1288 ();
 sg13g2_decap_8 FILLER_2_1295 ();
 sg13g2_decap_8 FILLER_2_1302 ();
 sg13g2_decap_4 FILLER_2_1309 ();
 sg13g2_fill_2 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_174 ();
 sg13g2_fill_1 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_fill_2 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_246 ();
 sg13g2_decap_4 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_4 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_fill_2 FILLER_3_339 ();
 sg13g2_fill_2 FILLER_3_367 ();
 sg13g2_fill_1 FILLER_3_369 ();
 sg13g2_decap_4 FILLER_3_377 ();
 sg13g2_decap_4 FILLER_3_385 ();
 sg13g2_fill_2 FILLER_3_389 ();
 sg13g2_fill_2 FILLER_3_422 ();
 sg13g2_decap_4 FILLER_3_476 ();
 sg13g2_fill_2 FILLER_3_480 ();
 sg13g2_fill_1 FILLER_3_534 ();
 sg13g2_decap_8 FILLER_3_549 ();
 sg13g2_fill_2 FILLER_3_556 ();
 sg13g2_fill_2 FILLER_3_576 ();
 sg13g2_fill_1 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_fill_1 FILLER_3_652 ();
 sg13g2_decap_8 FILLER_3_657 ();
 sg13g2_decap_4 FILLER_3_716 ();
 sg13g2_decap_4 FILLER_3_730 ();
 sg13g2_fill_1 FILLER_3_734 ();
 sg13g2_decap_4 FILLER_3_739 ();
 sg13g2_fill_1 FILLER_3_743 ();
 sg13g2_decap_4 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_820 ();
 sg13g2_fill_1 FILLER_3_827 ();
 sg13g2_decap_8 FILLER_3_895 ();
 sg13g2_fill_1 FILLER_3_902 ();
 sg13g2_fill_2 FILLER_3_913 ();
 sg13g2_decap_4 FILLER_3_934 ();
 sg13g2_fill_2 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_decap_8 FILLER_3_1026 ();
 sg13g2_decap_8 FILLER_3_1033 ();
 sg13g2_decap_8 FILLER_3_1040 ();
 sg13g2_decap_8 FILLER_3_1047 ();
 sg13g2_decap_8 FILLER_3_1054 ();
 sg13g2_decap_8 FILLER_3_1061 ();
 sg13g2_decap_8 FILLER_3_1068 ();
 sg13g2_decap_8 FILLER_3_1075 ();
 sg13g2_decap_8 FILLER_3_1082 ();
 sg13g2_decap_8 FILLER_3_1089 ();
 sg13g2_decap_8 FILLER_3_1096 ();
 sg13g2_decap_8 FILLER_3_1103 ();
 sg13g2_decap_8 FILLER_3_1110 ();
 sg13g2_decap_8 FILLER_3_1117 ();
 sg13g2_decap_8 FILLER_3_1124 ();
 sg13g2_decap_8 FILLER_3_1131 ();
 sg13g2_decap_8 FILLER_3_1138 ();
 sg13g2_decap_8 FILLER_3_1145 ();
 sg13g2_decap_8 FILLER_3_1152 ();
 sg13g2_decap_8 FILLER_3_1159 ();
 sg13g2_decap_8 FILLER_3_1166 ();
 sg13g2_decap_8 FILLER_3_1173 ();
 sg13g2_decap_8 FILLER_3_1180 ();
 sg13g2_decap_8 FILLER_3_1187 ();
 sg13g2_decap_8 FILLER_3_1194 ();
 sg13g2_decap_8 FILLER_3_1201 ();
 sg13g2_decap_8 FILLER_3_1208 ();
 sg13g2_decap_8 FILLER_3_1215 ();
 sg13g2_decap_8 FILLER_3_1222 ();
 sg13g2_decap_8 FILLER_3_1229 ();
 sg13g2_decap_8 FILLER_3_1236 ();
 sg13g2_decap_8 FILLER_3_1243 ();
 sg13g2_decap_8 FILLER_3_1250 ();
 sg13g2_decap_8 FILLER_3_1257 ();
 sg13g2_decap_8 FILLER_3_1264 ();
 sg13g2_decap_8 FILLER_3_1271 ();
 sg13g2_decap_8 FILLER_3_1278 ();
 sg13g2_decap_8 FILLER_3_1285 ();
 sg13g2_decap_8 FILLER_3_1292 ();
 sg13g2_decap_8 FILLER_3_1299 ();
 sg13g2_decap_8 FILLER_3_1306 ();
 sg13g2_fill_2 FILLER_3_1313 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_160 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_4 FILLER_4_179 ();
 sg13g2_fill_2 FILLER_4_183 ();
 sg13g2_fill_2 FILLER_4_229 ();
 sg13g2_fill_1 FILLER_4_231 ();
 sg13g2_decap_4 FILLER_4_258 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_269 ();
 sg13g2_fill_2 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_fill_2 FILLER_4_317 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_fill_2 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_450 ();
 sg13g2_decap_8 FILLER_4_457 ();
 sg13g2_fill_2 FILLER_4_464 ();
 sg13g2_fill_1 FILLER_4_466 ();
 sg13g2_decap_4 FILLER_4_477 ();
 sg13g2_decap_8 FILLER_4_491 ();
 sg13g2_fill_1 FILLER_4_498 ();
 sg13g2_decap_8 FILLER_4_503 ();
 sg13g2_fill_2 FILLER_4_519 ();
 sg13g2_decap_8 FILLER_4_598 ();
 sg13g2_decap_8 FILLER_4_605 ();
 sg13g2_fill_2 FILLER_4_612 ();
 sg13g2_decap_8 FILLER_4_628 ();
 sg13g2_decap_8 FILLER_4_635 ();
 sg13g2_decap_8 FILLER_4_668 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_fill_1 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_698 ();
 sg13g2_fill_2 FILLER_4_705 ();
 sg13g2_fill_1 FILLER_4_711 ();
 sg13g2_fill_2 FILLER_4_722 ();
 sg13g2_decap_8 FILLER_4_750 ();
 sg13g2_decap_4 FILLER_4_757 ();
 sg13g2_decap_8 FILLER_4_771 ();
 sg13g2_fill_2 FILLER_4_811 ();
 sg13g2_fill_1 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_fill_2 FILLER_4_847 ();
 sg13g2_decap_4 FILLER_4_879 ();
 sg13g2_fill_1 FILLER_4_883 ();
 sg13g2_fill_1 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_948 ();
 sg13g2_fill_1 FILLER_4_955 ();
 sg13g2_decap_8 FILLER_4_960 ();
 sg13g2_decap_4 FILLER_4_967 ();
 sg13g2_fill_1 FILLER_4_971 ();
 sg13g2_decap_8 FILLER_4_982 ();
 sg13g2_fill_1 FILLER_4_989 ();
 sg13g2_decap_8 FILLER_4_997 ();
 sg13g2_decap_8 FILLER_4_1004 ();
 sg13g2_decap_8 FILLER_4_1011 ();
 sg13g2_fill_1 FILLER_4_1018 ();
 sg13g2_decap_8 FILLER_4_1029 ();
 sg13g2_decap_8 FILLER_4_1036 ();
 sg13g2_decap_8 FILLER_4_1043 ();
 sg13g2_decap_8 FILLER_4_1050 ();
 sg13g2_decap_8 FILLER_4_1057 ();
 sg13g2_decap_8 FILLER_4_1064 ();
 sg13g2_decap_8 FILLER_4_1071 ();
 sg13g2_decap_8 FILLER_4_1078 ();
 sg13g2_decap_8 FILLER_4_1085 ();
 sg13g2_decap_8 FILLER_4_1092 ();
 sg13g2_decap_8 FILLER_4_1099 ();
 sg13g2_decap_8 FILLER_4_1106 ();
 sg13g2_decap_8 FILLER_4_1113 ();
 sg13g2_decap_8 FILLER_4_1120 ();
 sg13g2_decap_8 FILLER_4_1127 ();
 sg13g2_decap_8 FILLER_4_1134 ();
 sg13g2_decap_8 FILLER_4_1141 ();
 sg13g2_decap_8 FILLER_4_1148 ();
 sg13g2_decap_8 FILLER_4_1155 ();
 sg13g2_decap_8 FILLER_4_1162 ();
 sg13g2_decap_8 FILLER_4_1169 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_decap_8 FILLER_4_1183 ();
 sg13g2_decap_8 FILLER_4_1190 ();
 sg13g2_decap_8 FILLER_4_1197 ();
 sg13g2_decap_8 FILLER_4_1204 ();
 sg13g2_decap_8 FILLER_4_1211 ();
 sg13g2_decap_8 FILLER_4_1218 ();
 sg13g2_decap_8 FILLER_4_1225 ();
 sg13g2_decap_8 FILLER_4_1232 ();
 sg13g2_decap_8 FILLER_4_1239 ();
 sg13g2_decap_8 FILLER_4_1246 ();
 sg13g2_decap_8 FILLER_4_1253 ();
 sg13g2_decap_8 FILLER_4_1260 ();
 sg13g2_decap_8 FILLER_4_1267 ();
 sg13g2_decap_8 FILLER_4_1274 ();
 sg13g2_decap_8 FILLER_4_1281 ();
 sg13g2_decap_8 FILLER_4_1288 ();
 sg13g2_decap_8 FILLER_4_1295 ();
 sg13g2_decap_8 FILLER_4_1302 ();
 sg13g2_decap_4 FILLER_4_1309 ();
 sg13g2_fill_2 FILLER_4_1313 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_156 ();
 sg13g2_fill_2 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_decap_4 FILLER_5_201 ();
 sg13g2_decap_4 FILLER_5_209 ();
 sg13g2_decap_4 FILLER_5_218 ();
 sg13g2_fill_2 FILLER_5_222 ();
 sg13g2_fill_2 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_4 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_264 ();
 sg13g2_fill_1 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_287 ();
 sg13g2_decap_4 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_345 ();
 sg13g2_fill_1 FILLER_5_370 ();
 sg13g2_fill_1 FILLER_5_390 ();
 sg13g2_fill_2 FILLER_5_402 ();
 sg13g2_fill_1 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_418 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_fill_2 FILLER_5_480 ();
 sg13g2_fill_2 FILLER_5_496 ();
 sg13g2_fill_1 FILLER_5_498 ();
 sg13g2_decap_8 FILLER_5_528 ();
 sg13g2_fill_2 FILLER_5_535 ();
 sg13g2_fill_1 FILLER_5_537 ();
 sg13g2_decap_8 FILLER_5_548 ();
 sg13g2_decap_4 FILLER_5_555 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_fill_1 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_593 ();
 sg13g2_decap_4 FILLER_5_600 ();
 sg13g2_fill_1 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_631 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_fill_2 FILLER_5_645 ();
 sg13g2_fill_1 FILLER_5_657 ();
 sg13g2_decap_8 FILLER_5_673 ();
 sg13g2_fill_1 FILLER_5_680 ();
 sg13g2_fill_1 FILLER_5_695 ();
 sg13g2_fill_2 FILLER_5_722 ();
 sg13g2_fill_1 FILLER_5_724 ();
 sg13g2_fill_2 FILLER_5_735 ();
 sg13g2_decap_4 FILLER_5_741 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_decap_8 FILLER_5_778 ();
 sg13g2_fill_1 FILLER_5_785 ();
 sg13g2_fill_2 FILLER_5_790 ();
 sg13g2_decap_4 FILLER_5_796 ();
 sg13g2_fill_1 FILLER_5_810 ();
 sg13g2_decap_4 FILLER_5_821 ();
 sg13g2_fill_1 FILLER_5_829 ();
 sg13g2_decap_4 FILLER_5_866 ();
 sg13g2_fill_1 FILLER_5_870 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_fill_2 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_899 ();
 sg13g2_decap_8 FILLER_5_906 ();
 sg13g2_fill_2 FILLER_5_913 ();
 sg13g2_decap_4 FILLER_5_925 ();
 sg13g2_fill_2 FILLER_5_933 ();
 sg13g2_decap_8 FILLER_5_971 ();
 sg13g2_fill_2 FILLER_5_978 ();
 sg13g2_decap_8 FILLER_5_1058 ();
 sg13g2_decap_8 FILLER_5_1065 ();
 sg13g2_decap_8 FILLER_5_1072 ();
 sg13g2_decap_8 FILLER_5_1079 ();
 sg13g2_decap_8 FILLER_5_1086 ();
 sg13g2_decap_8 FILLER_5_1093 ();
 sg13g2_decap_8 FILLER_5_1100 ();
 sg13g2_decap_8 FILLER_5_1107 ();
 sg13g2_decap_8 FILLER_5_1114 ();
 sg13g2_decap_8 FILLER_5_1121 ();
 sg13g2_decap_8 FILLER_5_1128 ();
 sg13g2_decap_8 FILLER_5_1135 ();
 sg13g2_decap_8 FILLER_5_1142 ();
 sg13g2_decap_8 FILLER_5_1149 ();
 sg13g2_decap_8 FILLER_5_1156 ();
 sg13g2_decap_8 FILLER_5_1163 ();
 sg13g2_decap_8 FILLER_5_1170 ();
 sg13g2_decap_8 FILLER_5_1177 ();
 sg13g2_decap_8 FILLER_5_1184 ();
 sg13g2_decap_8 FILLER_5_1191 ();
 sg13g2_decap_8 FILLER_5_1198 ();
 sg13g2_decap_8 FILLER_5_1205 ();
 sg13g2_decap_8 FILLER_5_1212 ();
 sg13g2_decap_8 FILLER_5_1219 ();
 sg13g2_decap_8 FILLER_5_1226 ();
 sg13g2_decap_8 FILLER_5_1233 ();
 sg13g2_decap_8 FILLER_5_1240 ();
 sg13g2_decap_8 FILLER_5_1247 ();
 sg13g2_decap_8 FILLER_5_1254 ();
 sg13g2_decap_8 FILLER_5_1261 ();
 sg13g2_decap_8 FILLER_5_1268 ();
 sg13g2_decap_8 FILLER_5_1275 ();
 sg13g2_decap_8 FILLER_5_1282 ();
 sg13g2_decap_8 FILLER_5_1289 ();
 sg13g2_decap_8 FILLER_5_1296 ();
 sg13g2_decap_8 FILLER_5_1303 ();
 sg13g2_decap_4 FILLER_5_1310 ();
 sg13g2_fill_1 FILLER_5_1314 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_decap_4 FILLER_6_205 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_fill_1 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_fill_2 FILLER_6_325 ();
 sg13g2_fill_2 FILLER_6_334 ();
 sg13g2_decap_4 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_344 ();
 sg13g2_fill_2 FILLER_6_371 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_2 FILLER_6_383 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_fill_1 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_435 ();
 sg13g2_fill_2 FILLER_6_453 ();
 sg13g2_fill_1 FILLER_6_455 ();
 sg13g2_fill_2 FILLER_6_474 ();
 sg13g2_fill_1 FILLER_6_476 ();
 sg13g2_fill_2 FILLER_6_490 ();
 sg13g2_fill_1 FILLER_6_498 ();
 sg13g2_fill_1 FILLER_6_511 ();
 sg13g2_fill_2 FILLER_6_523 ();
 sg13g2_decap_8 FILLER_6_533 ();
 sg13g2_decap_8 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_decap_8 FILLER_6_580 ();
 sg13g2_fill_2 FILLER_6_587 ();
 sg13g2_decap_4 FILLER_6_610 ();
 sg13g2_fill_1 FILLER_6_614 ();
 sg13g2_decap_4 FILLER_6_619 ();
 sg13g2_fill_2 FILLER_6_710 ();
 sg13g2_decap_4 FILLER_6_722 ();
 sg13g2_fill_1 FILLER_6_755 ();
 sg13g2_decap_4 FILLER_6_760 ();
 sg13g2_fill_1 FILLER_6_764 ();
 sg13g2_decap_4 FILLER_6_811 ();
 sg13g2_fill_1 FILLER_6_815 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_4 FILLER_6_847 ();
 sg13g2_decap_4 FILLER_6_855 ();
 sg13g2_fill_1 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_874 ();
 sg13g2_decap_8 FILLER_6_881 ();
 sg13g2_fill_1 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_910 ();
 sg13g2_fill_1 FILLER_6_917 ();
 sg13g2_fill_2 FILLER_6_944 ();
 sg13g2_fill_2 FILLER_6_956 ();
 sg13g2_fill_1 FILLER_6_958 ();
 sg13g2_decap_4 FILLER_6_983 ();
 sg13g2_fill_2 FILLER_6_987 ();
 sg13g2_fill_1 FILLER_6_1009 ();
 sg13g2_fill_2 FILLER_6_1024 ();
 sg13g2_fill_1 FILLER_6_1026 ();
 sg13g2_decap_4 FILLER_6_1037 ();
 sg13g2_fill_1 FILLER_6_1041 ();
 sg13g2_decap_8 FILLER_6_1046 ();
 sg13g2_decap_8 FILLER_6_1053 ();
 sg13g2_decap_8 FILLER_6_1060 ();
 sg13g2_decap_8 FILLER_6_1067 ();
 sg13g2_decap_8 FILLER_6_1074 ();
 sg13g2_decap_8 FILLER_6_1081 ();
 sg13g2_decap_8 FILLER_6_1088 ();
 sg13g2_decap_8 FILLER_6_1095 ();
 sg13g2_decap_8 FILLER_6_1102 ();
 sg13g2_decap_8 FILLER_6_1109 ();
 sg13g2_decap_8 FILLER_6_1116 ();
 sg13g2_decap_8 FILLER_6_1123 ();
 sg13g2_decap_8 FILLER_6_1130 ();
 sg13g2_decap_8 FILLER_6_1137 ();
 sg13g2_decap_8 FILLER_6_1144 ();
 sg13g2_decap_8 FILLER_6_1151 ();
 sg13g2_decap_8 FILLER_6_1158 ();
 sg13g2_decap_8 FILLER_6_1165 ();
 sg13g2_decap_8 FILLER_6_1172 ();
 sg13g2_decap_8 FILLER_6_1179 ();
 sg13g2_decap_8 FILLER_6_1186 ();
 sg13g2_decap_8 FILLER_6_1193 ();
 sg13g2_decap_8 FILLER_6_1200 ();
 sg13g2_decap_8 FILLER_6_1207 ();
 sg13g2_decap_8 FILLER_6_1214 ();
 sg13g2_decap_8 FILLER_6_1221 ();
 sg13g2_decap_8 FILLER_6_1228 ();
 sg13g2_decap_8 FILLER_6_1235 ();
 sg13g2_decap_8 FILLER_6_1242 ();
 sg13g2_decap_8 FILLER_6_1249 ();
 sg13g2_decap_8 FILLER_6_1256 ();
 sg13g2_decap_8 FILLER_6_1263 ();
 sg13g2_decap_8 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1277 ();
 sg13g2_decap_8 FILLER_6_1284 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_fill_2 FILLER_6_1312 ();
 sg13g2_fill_1 FILLER_6_1314 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_1 FILLER_7_98 ();
 sg13g2_decap_4 FILLER_7_125 ();
 sg13g2_fill_1 FILLER_7_129 ();
 sg13g2_decap_8 FILLER_7_134 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_decap_4 FILLER_7_148 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_decap_4 FILLER_7_176 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_2 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_decap_4 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_2 FILLER_7_323 ();
 sg13g2_decap_4 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_4 FILLER_7_417 ();
 sg13g2_fill_2 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_7_431 ();
 sg13g2_fill_2 FILLER_7_461 ();
 sg13g2_fill_1 FILLER_7_463 ();
 sg13g2_fill_2 FILLER_7_479 ();
 sg13g2_decap_4 FILLER_7_496 ();
 sg13g2_fill_1 FILLER_7_500 ();
 sg13g2_fill_1 FILLER_7_514 ();
 sg13g2_decap_4 FILLER_7_539 ();
 sg13g2_fill_2 FILLER_7_543 ();
 sg13g2_decap_4 FILLER_7_585 ();
 sg13g2_fill_2 FILLER_7_610 ();
 sg13g2_fill_1 FILLER_7_612 ();
 sg13g2_fill_2 FILLER_7_644 ();
 sg13g2_fill_2 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_666 ();
 sg13g2_decap_4 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_677 ();
 sg13g2_decap_4 FILLER_7_689 ();
 sg13g2_fill_2 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_731 ();
 sg13g2_decap_8 FILLER_7_738 ();
 sg13g2_decap_8 FILLER_7_745 ();
 sg13g2_decap_8 FILLER_7_773 ();
 sg13g2_decap_4 FILLER_7_780 ();
 sg13g2_fill_2 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_4 FILLER_7_804 ();
 sg13g2_decap_4 FILLER_7_813 ();
 sg13g2_fill_1 FILLER_7_817 ();
 sg13g2_decap_4 FILLER_7_823 ();
 sg13g2_decap_8 FILLER_7_837 ();
 sg13g2_decap_8 FILLER_7_844 ();
 sg13g2_decap_4 FILLER_7_851 ();
 sg13g2_fill_1 FILLER_7_855 ();
 sg13g2_fill_2 FILLER_7_874 ();
 sg13g2_fill_1 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_900 ();
 sg13g2_decap_8 FILLER_7_907 ();
 sg13g2_decap_8 FILLER_7_914 ();
 sg13g2_fill_2 FILLER_7_957 ();
 sg13g2_decap_4 FILLER_7_979 ();
 sg13g2_fill_2 FILLER_7_983 ();
 sg13g2_fill_2 FILLER_7_995 ();
 sg13g2_fill_1 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1024 ();
 sg13g2_decap_8 FILLER_7_1045 ();
 sg13g2_decap_8 FILLER_7_1056 ();
 sg13g2_decap_8 FILLER_7_1063 ();
 sg13g2_decap_8 FILLER_7_1070 ();
 sg13g2_decap_8 FILLER_7_1077 ();
 sg13g2_decap_8 FILLER_7_1084 ();
 sg13g2_decap_8 FILLER_7_1091 ();
 sg13g2_decap_8 FILLER_7_1098 ();
 sg13g2_decap_8 FILLER_7_1105 ();
 sg13g2_decap_8 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1119 ();
 sg13g2_decap_8 FILLER_7_1126 ();
 sg13g2_decap_8 FILLER_7_1133 ();
 sg13g2_decap_8 FILLER_7_1140 ();
 sg13g2_decap_8 FILLER_7_1147 ();
 sg13g2_decap_8 FILLER_7_1154 ();
 sg13g2_decap_8 FILLER_7_1161 ();
 sg13g2_decap_8 FILLER_7_1168 ();
 sg13g2_decap_8 FILLER_7_1175 ();
 sg13g2_decap_8 FILLER_7_1182 ();
 sg13g2_decap_8 FILLER_7_1189 ();
 sg13g2_decap_8 FILLER_7_1196 ();
 sg13g2_decap_8 FILLER_7_1203 ();
 sg13g2_decap_8 FILLER_7_1210 ();
 sg13g2_decap_8 FILLER_7_1217 ();
 sg13g2_decap_8 FILLER_7_1224 ();
 sg13g2_decap_8 FILLER_7_1231 ();
 sg13g2_decap_8 FILLER_7_1238 ();
 sg13g2_decap_8 FILLER_7_1245 ();
 sg13g2_decap_8 FILLER_7_1252 ();
 sg13g2_decap_8 FILLER_7_1259 ();
 sg13g2_decap_8 FILLER_7_1266 ();
 sg13g2_decap_8 FILLER_7_1273 ();
 sg13g2_decap_8 FILLER_7_1280 ();
 sg13g2_decap_8 FILLER_7_1287 ();
 sg13g2_decap_8 FILLER_7_1294 ();
 sg13g2_decap_8 FILLER_7_1301 ();
 sg13g2_decap_8 FILLER_7_1308 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_4 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_decap_4 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_299 ();
 sg13g2_decap_4 FILLER_8_313 ();
 sg13g2_decap_4 FILLER_8_324 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_4 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_fill_2 FILLER_8_421 ();
 sg13g2_fill_2 FILLER_8_440 ();
 sg13g2_fill_1 FILLER_8_442 ();
 sg13g2_fill_2 FILLER_8_449 ();
 sg13g2_fill_2 FILLER_8_471 ();
 sg13g2_fill_1 FILLER_8_473 ();
 sg13g2_fill_1 FILLER_8_493 ();
 sg13g2_decap_4 FILLER_8_505 ();
 sg13g2_decap_8 FILLER_8_535 ();
 sg13g2_decap_8 FILLER_8_542 ();
 sg13g2_decap_4 FILLER_8_549 ();
 sg13g2_fill_2 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_559 ();
 sg13g2_fill_2 FILLER_8_566 ();
 sg13g2_fill_1 FILLER_8_568 ();
 sg13g2_fill_2 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_596 ();
 sg13g2_fill_2 FILLER_8_633 ();
 sg13g2_fill_2 FILLER_8_661 ();
 sg13g2_decap_4 FILLER_8_689 ();
 sg13g2_fill_2 FILLER_8_719 ();
 sg13g2_fill_1 FILLER_8_721 ();
 sg13g2_fill_2 FILLER_8_802 ();
 sg13g2_fill_1 FILLER_8_804 ();
 sg13g2_fill_1 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_fill_1 FILLER_8_878 ();
 sg13g2_fill_2 FILLER_8_930 ();
 sg13g2_decap_8 FILLER_8_936 ();
 sg13g2_decap_4 FILLER_8_943 ();
 sg13g2_fill_2 FILLER_8_947 ();
 sg13g2_fill_1 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_fill_1 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_1072 ();
 sg13g2_decap_8 FILLER_8_1079 ();
 sg13g2_decap_8 FILLER_8_1086 ();
 sg13g2_decap_8 FILLER_8_1093 ();
 sg13g2_decap_8 FILLER_8_1100 ();
 sg13g2_decap_8 FILLER_8_1107 ();
 sg13g2_decap_8 FILLER_8_1114 ();
 sg13g2_decap_8 FILLER_8_1121 ();
 sg13g2_decap_8 FILLER_8_1128 ();
 sg13g2_decap_8 FILLER_8_1135 ();
 sg13g2_decap_8 FILLER_8_1142 ();
 sg13g2_decap_8 FILLER_8_1149 ();
 sg13g2_decap_8 FILLER_8_1156 ();
 sg13g2_decap_8 FILLER_8_1163 ();
 sg13g2_decap_8 FILLER_8_1170 ();
 sg13g2_decap_8 FILLER_8_1177 ();
 sg13g2_decap_8 FILLER_8_1184 ();
 sg13g2_decap_8 FILLER_8_1191 ();
 sg13g2_decap_8 FILLER_8_1198 ();
 sg13g2_decap_8 FILLER_8_1205 ();
 sg13g2_decap_8 FILLER_8_1212 ();
 sg13g2_decap_8 FILLER_8_1219 ();
 sg13g2_decap_8 FILLER_8_1226 ();
 sg13g2_decap_8 FILLER_8_1233 ();
 sg13g2_decap_8 FILLER_8_1240 ();
 sg13g2_decap_8 FILLER_8_1247 ();
 sg13g2_decap_8 FILLER_8_1254 ();
 sg13g2_decap_8 FILLER_8_1261 ();
 sg13g2_decap_8 FILLER_8_1268 ();
 sg13g2_decap_8 FILLER_8_1275 ();
 sg13g2_decap_8 FILLER_8_1282 ();
 sg13g2_decap_8 FILLER_8_1289 ();
 sg13g2_decap_8 FILLER_8_1296 ();
 sg13g2_decap_8 FILLER_8_1303 ();
 sg13g2_decap_4 FILLER_8_1310 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_26 ();
 sg13g2_decap_8 FILLER_9_33 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_decap_4 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_52 ();
 sg13g2_decap_4 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_61 ();
 sg13g2_decap_8 FILLER_9_65 ();
 sg13g2_decap_8 FILLER_9_72 ();
 sg13g2_decap_4 FILLER_9_79 ();
 sg13g2_fill_2 FILLER_9_83 ();
 sg13g2_fill_2 FILLER_9_111 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_4 FILLER_9_175 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_4 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_387 ();
 sg13g2_decap_4 FILLER_9_394 ();
 sg13g2_fill_2 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_fill_2 FILLER_9_416 ();
 sg13g2_decap_4 FILLER_9_423 ();
 sg13g2_decap_8 FILLER_9_435 ();
 sg13g2_decap_4 FILLER_9_442 ();
 sg13g2_fill_1 FILLER_9_446 ();
 sg13g2_decap_8 FILLER_9_457 ();
 sg13g2_fill_2 FILLER_9_464 ();
 sg13g2_fill_1 FILLER_9_466 ();
 sg13g2_fill_2 FILLER_9_477 ();
 sg13g2_fill_1 FILLER_9_479 ();
 sg13g2_decap_8 FILLER_9_485 ();
 sg13g2_fill_2 FILLER_9_492 ();
 sg13g2_decap_4 FILLER_9_514 ();
 sg13g2_fill_2 FILLER_9_518 ();
 sg13g2_decap_4 FILLER_9_525 ();
 sg13g2_fill_1 FILLER_9_533 ();
 sg13g2_decap_4 FILLER_9_570 ();
 sg13g2_fill_1 FILLER_9_574 ();
 sg13g2_fill_2 FILLER_9_596 ();
 sg13g2_fill_2 FILLER_9_634 ();
 sg13g2_fill_1 FILLER_9_636 ();
 sg13g2_fill_1 FILLER_9_647 ();
 sg13g2_decap_4 FILLER_9_669 ();
 sg13g2_fill_1 FILLER_9_673 ();
 sg13g2_fill_2 FILLER_9_678 ();
 sg13g2_decap_4 FILLER_9_690 ();
 sg13g2_fill_1 FILLER_9_694 ();
 sg13g2_decap_8 FILLER_9_720 ();
 sg13g2_decap_8 FILLER_9_741 ();
 sg13g2_decap_4 FILLER_9_768 ();
 sg13g2_fill_1 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_fill_2 FILLER_9_833 ();
 sg13g2_fill_1 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_fill_1 FILLER_9_851 ();
 sg13g2_fill_1 FILLER_9_864 ();
 sg13g2_fill_1 FILLER_9_883 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_fill_1 FILLER_9_900 ();
 sg13g2_fill_2 FILLER_9_909 ();
 sg13g2_fill_2 FILLER_9_965 ();
 sg13g2_decap_8 FILLER_9_972 ();
 sg13g2_fill_2 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_1004 ();
 sg13g2_fill_2 FILLER_9_1011 ();
 sg13g2_decap_8 FILLER_9_1023 ();
 sg13g2_decap_4 FILLER_9_1030 ();
 sg13g2_fill_2 FILLER_9_1034 ();
 sg13g2_decap_8 FILLER_9_1041 ();
 sg13g2_fill_2 FILLER_9_1048 ();
 sg13g2_decap_8 FILLER_9_1086 ();
 sg13g2_decap_8 FILLER_9_1093 ();
 sg13g2_decap_8 FILLER_9_1100 ();
 sg13g2_decap_8 FILLER_9_1107 ();
 sg13g2_decap_8 FILLER_9_1114 ();
 sg13g2_decap_8 FILLER_9_1121 ();
 sg13g2_decap_8 FILLER_9_1128 ();
 sg13g2_decap_8 FILLER_9_1135 ();
 sg13g2_decap_8 FILLER_9_1142 ();
 sg13g2_decap_8 FILLER_9_1149 ();
 sg13g2_decap_8 FILLER_9_1156 ();
 sg13g2_decap_8 FILLER_9_1163 ();
 sg13g2_decap_8 FILLER_9_1170 ();
 sg13g2_decap_8 FILLER_9_1177 ();
 sg13g2_decap_8 FILLER_9_1184 ();
 sg13g2_decap_8 FILLER_9_1191 ();
 sg13g2_decap_8 FILLER_9_1198 ();
 sg13g2_decap_8 FILLER_9_1205 ();
 sg13g2_decap_8 FILLER_9_1212 ();
 sg13g2_decap_8 FILLER_9_1219 ();
 sg13g2_decap_8 FILLER_9_1226 ();
 sg13g2_decap_8 FILLER_9_1233 ();
 sg13g2_decap_8 FILLER_9_1240 ();
 sg13g2_decap_8 FILLER_9_1247 ();
 sg13g2_decap_8 FILLER_9_1254 ();
 sg13g2_decap_8 FILLER_9_1261 ();
 sg13g2_decap_8 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1275 ();
 sg13g2_decap_8 FILLER_9_1282 ();
 sg13g2_decap_8 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1296 ();
 sg13g2_decap_8 FILLER_9_1303 ();
 sg13g2_decap_4 FILLER_9_1310 ();
 sg13g2_fill_1 FILLER_9_1314 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_68 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_4 FILLER_10_81 ();
 sg13g2_fill_1 FILLER_10_85 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_decap_4 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_139 ();
 sg13g2_fill_2 FILLER_10_150 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_2 FILLER_10_258 ();
 sg13g2_fill_1 FILLER_10_260 ();
 sg13g2_fill_1 FILLER_10_270 ();
 sg13g2_fill_1 FILLER_10_296 ();
 sg13g2_decap_4 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_decap_4 FILLER_10_320 ();
 sg13g2_fill_2 FILLER_10_335 ();
 sg13g2_fill_2 FILLER_10_341 ();
 sg13g2_decap_4 FILLER_10_352 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_fill_2 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_386 ();
 sg13g2_decap_4 FILLER_10_413 ();
 sg13g2_fill_2 FILLER_10_462 ();
 sg13g2_fill_1 FILLER_10_464 ();
 sg13g2_decap_4 FILLER_10_483 ();
 sg13g2_decap_4 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_545 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_fill_1 FILLER_10_592 ();
 sg13g2_decap_4 FILLER_10_603 ();
 sg13g2_fill_1 FILLER_10_607 ();
 sg13g2_decap_4 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_652 ();
 sg13g2_decap_4 FILLER_10_659 ();
 sg13g2_fill_1 FILLER_10_663 ();
 sg13g2_decap_4 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_715 ();
 sg13g2_decap_4 FILLER_10_751 ();
 sg13g2_fill_2 FILLER_10_755 ();
 sg13g2_fill_1 FILLER_10_765 ();
 sg13g2_fill_1 FILLER_10_776 ();
 sg13g2_decap_4 FILLER_10_781 ();
 sg13g2_fill_1 FILLER_10_785 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_4 FILLER_10_802 ();
 sg13g2_fill_2 FILLER_10_816 ();
 sg13g2_fill_1 FILLER_10_823 ();
 sg13g2_fill_1 FILLER_10_864 ();
 sg13g2_fill_2 FILLER_10_878 ();
 sg13g2_fill_2 FILLER_10_916 ();
 sg13g2_decap_8 FILLER_10_926 ();
 sg13g2_decap_4 FILLER_10_937 ();
 sg13g2_fill_2 FILLER_10_941 ();
 sg13g2_fill_2 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_972 ();
 sg13g2_fill_1 FILLER_10_979 ();
 sg13g2_decap_4 FILLER_10_983 ();
 sg13g2_fill_2 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_999 ();
 sg13g2_fill_2 FILLER_10_1016 ();
 sg13g2_fill_1 FILLER_10_1070 ();
 sg13g2_decap_4 FILLER_10_1075 ();
 sg13g2_fill_2 FILLER_10_1083 ();
 sg13g2_decap_8 FILLER_10_1095 ();
 sg13g2_decap_8 FILLER_10_1102 ();
 sg13g2_decap_8 FILLER_10_1109 ();
 sg13g2_decap_8 FILLER_10_1116 ();
 sg13g2_decap_8 FILLER_10_1123 ();
 sg13g2_decap_8 FILLER_10_1130 ();
 sg13g2_decap_8 FILLER_10_1137 ();
 sg13g2_decap_8 FILLER_10_1144 ();
 sg13g2_decap_8 FILLER_10_1151 ();
 sg13g2_decap_8 FILLER_10_1158 ();
 sg13g2_decap_8 FILLER_10_1165 ();
 sg13g2_decap_8 FILLER_10_1172 ();
 sg13g2_decap_8 FILLER_10_1179 ();
 sg13g2_decap_8 FILLER_10_1186 ();
 sg13g2_decap_8 FILLER_10_1193 ();
 sg13g2_decap_8 FILLER_10_1200 ();
 sg13g2_decap_8 FILLER_10_1207 ();
 sg13g2_decap_8 FILLER_10_1214 ();
 sg13g2_decap_8 FILLER_10_1221 ();
 sg13g2_decap_8 FILLER_10_1228 ();
 sg13g2_decap_8 FILLER_10_1235 ();
 sg13g2_decap_8 FILLER_10_1242 ();
 sg13g2_decap_8 FILLER_10_1249 ();
 sg13g2_decap_8 FILLER_10_1256 ();
 sg13g2_decap_8 FILLER_10_1263 ();
 sg13g2_decap_8 FILLER_10_1270 ();
 sg13g2_decap_8 FILLER_10_1277 ();
 sg13g2_decap_8 FILLER_10_1284 ();
 sg13g2_decap_8 FILLER_10_1291 ();
 sg13g2_decap_8 FILLER_10_1298 ();
 sg13g2_decap_8 FILLER_10_1305 ();
 sg13g2_fill_2 FILLER_10_1312 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_32 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_2 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_1 FILLER_11_333 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_373 ();
 sg13g2_fill_1 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_fill_1 FILLER_11_410 ();
 sg13g2_fill_2 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_430 ();
 sg13g2_decap_4 FILLER_11_437 ();
 sg13g2_fill_1 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_464 ();
 sg13g2_decap_8 FILLER_11_471 ();
 sg13g2_fill_1 FILLER_11_483 ();
 sg13g2_fill_1 FILLER_11_497 ();
 sg13g2_fill_1 FILLER_11_502 ();
 sg13g2_fill_2 FILLER_11_511 ();
 sg13g2_fill_2 FILLER_11_561 ();
 sg13g2_fill_1 FILLER_11_571 ();
 sg13g2_decap_4 FILLER_11_632 ();
 sg13g2_fill_2 FILLER_11_648 ();
 sg13g2_fill_2 FILLER_11_671 ();
 sg13g2_decap_8 FILLER_11_685 ();
 sg13g2_decap_8 FILLER_11_692 ();
 sg13g2_decap_8 FILLER_11_699 ();
 sg13g2_fill_2 FILLER_11_706 ();
 sg13g2_fill_1 FILLER_11_708 ();
 sg13g2_decap_8 FILLER_11_717 ();
 sg13g2_fill_1 FILLER_11_724 ();
 sg13g2_fill_2 FILLER_11_737 ();
 sg13g2_fill_2 FILLER_11_754 ();
 sg13g2_fill_1 FILLER_11_792 ();
 sg13g2_decap_4 FILLER_11_811 ();
 sg13g2_fill_2 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_4 FILLER_11_842 ();
 sg13g2_fill_2 FILLER_11_846 ();
 sg13g2_decap_8 FILLER_11_852 ();
 sg13g2_fill_2 FILLER_11_867 ();
 sg13g2_fill_1 FILLER_11_869 ();
 sg13g2_fill_2 FILLER_11_875 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_4 FILLER_11_893 ();
 sg13g2_fill_2 FILLER_11_901 ();
 sg13g2_fill_1 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_909 ();
 sg13g2_fill_2 FILLER_11_916 ();
 sg13g2_fill_2 FILLER_11_936 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_fill_1 FILLER_11_949 ();
 sg13g2_fill_2 FILLER_11_955 ();
 sg13g2_fill_1 FILLER_11_993 ();
 sg13g2_decap_8 FILLER_11_1020 ();
 sg13g2_fill_2 FILLER_11_1027 ();
 sg13g2_fill_1 FILLER_11_1033 ();
 sg13g2_decap_8 FILLER_11_1058 ();
 sg13g2_decap_4 FILLER_11_1065 ();
 sg13g2_decap_8 FILLER_11_1095 ();
 sg13g2_decap_8 FILLER_11_1102 ();
 sg13g2_decap_8 FILLER_11_1109 ();
 sg13g2_decap_8 FILLER_11_1116 ();
 sg13g2_decap_8 FILLER_11_1123 ();
 sg13g2_decap_8 FILLER_11_1130 ();
 sg13g2_decap_8 FILLER_11_1137 ();
 sg13g2_decap_8 FILLER_11_1144 ();
 sg13g2_decap_8 FILLER_11_1151 ();
 sg13g2_decap_8 FILLER_11_1158 ();
 sg13g2_decap_8 FILLER_11_1165 ();
 sg13g2_decap_8 FILLER_11_1172 ();
 sg13g2_decap_8 FILLER_11_1179 ();
 sg13g2_decap_8 FILLER_11_1186 ();
 sg13g2_decap_8 FILLER_11_1193 ();
 sg13g2_decap_8 FILLER_11_1200 ();
 sg13g2_decap_8 FILLER_11_1207 ();
 sg13g2_decap_8 FILLER_11_1214 ();
 sg13g2_decap_8 FILLER_11_1221 ();
 sg13g2_decap_8 FILLER_11_1228 ();
 sg13g2_decap_8 FILLER_11_1235 ();
 sg13g2_decap_8 FILLER_11_1242 ();
 sg13g2_decap_8 FILLER_11_1249 ();
 sg13g2_decap_8 FILLER_11_1256 ();
 sg13g2_decap_8 FILLER_11_1263 ();
 sg13g2_decap_8 FILLER_11_1270 ();
 sg13g2_decap_8 FILLER_11_1277 ();
 sg13g2_decap_8 FILLER_11_1284 ();
 sg13g2_decap_8 FILLER_11_1291 ();
 sg13g2_decap_8 FILLER_11_1298 ();
 sg13g2_decap_8 FILLER_11_1305 ();
 sg13g2_fill_2 FILLER_11_1312 ();
 sg13g2_fill_1 FILLER_11_1314 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_decap_4 FILLER_12_9 ();
 sg13g2_fill_1 FILLER_12_13 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_2 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_decap_8 FILLER_12_99 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_fill_2 FILLER_12_138 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_decap_4 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_2 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_244 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_310 ();
 sg13g2_fill_1 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_4 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_decap_4 FILLER_12_416 ();
 sg13g2_fill_1 FILLER_12_420 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_2 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_12_447 ();
 sg13g2_decap_4 FILLER_12_471 ();
 sg13g2_decap_4 FILLER_12_482 ();
 sg13g2_decap_4 FILLER_12_491 ();
 sg13g2_fill_1 FILLER_12_495 ();
 sg13g2_decap_8 FILLER_12_527 ();
 sg13g2_fill_1 FILLER_12_534 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_4 FILLER_12_546 ();
 sg13g2_fill_2 FILLER_12_550 ();
 sg13g2_fill_1 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_4 FILLER_12_613 ();
 sg13g2_fill_2 FILLER_12_617 ();
 sg13g2_decap_8 FILLER_12_632 ();
 sg13g2_decap_4 FILLER_12_639 ();
 sg13g2_fill_2 FILLER_12_643 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_4 FILLER_12_670 ();
 sg13g2_fill_2 FILLER_12_674 ();
 sg13g2_fill_1 FILLER_12_682 ();
 sg13g2_fill_2 FILLER_12_692 ();
 sg13g2_fill_1 FILLER_12_694 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_fill_2 FILLER_12_707 ();
 sg13g2_fill_2 FILLER_12_732 ();
 sg13g2_fill_1 FILLER_12_734 ();
 sg13g2_decap_8 FILLER_12_751 ();
 sg13g2_decap_8 FILLER_12_758 ();
 sg13g2_decap_4 FILLER_12_765 ();
 sg13g2_decap_4 FILLER_12_779 ();
 sg13g2_fill_1 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_787 ();
 sg13g2_decap_4 FILLER_12_794 ();
 sg13g2_fill_2 FILLER_12_798 ();
 sg13g2_decap_4 FILLER_12_814 ();
 sg13g2_fill_1 FILLER_12_818 ();
 sg13g2_fill_1 FILLER_12_868 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_fill_2 FILLER_12_977 ();
 sg13g2_fill_1 FILLER_12_1049 ();
 sg13g2_decap_8 FILLER_12_1120 ();
 sg13g2_decap_8 FILLER_12_1127 ();
 sg13g2_decap_8 FILLER_12_1134 ();
 sg13g2_decap_8 FILLER_12_1141 ();
 sg13g2_decap_8 FILLER_12_1148 ();
 sg13g2_decap_8 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1169 ();
 sg13g2_decap_8 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1190 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_decap_8 FILLER_12_1204 ();
 sg13g2_decap_8 FILLER_12_1211 ();
 sg13g2_decap_8 FILLER_12_1218 ();
 sg13g2_decap_8 FILLER_12_1225 ();
 sg13g2_decap_8 FILLER_12_1232 ();
 sg13g2_decap_8 FILLER_12_1239 ();
 sg13g2_decap_8 FILLER_12_1246 ();
 sg13g2_decap_8 FILLER_12_1253 ();
 sg13g2_decap_8 FILLER_12_1260 ();
 sg13g2_decap_8 FILLER_12_1267 ();
 sg13g2_decap_8 FILLER_12_1274 ();
 sg13g2_decap_8 FILLER_12_1281 ();
 sg13g2_decap_8 FILLER_12_1288 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_4 FILLER_12_1309 ();
 sg13g2_fill_2 FILLER_12_1313 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_decap_4 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_fill_2 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_2 FILLER_13_94 ();
 sg13g2_fill_2 FILLER_13_100 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_decap_4 FILLER_13_108 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_301 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_fill_2 FILLER_13_356 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_decap_4 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_13_443 ();
 sg13g2_fill_1 FILLER_13_455 ();
 sg13g2_fill_2 FILLER_13_465 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_482 ();
 sg13g2_decap_8 FILLER_13_496 ();
 sg13g2_fill_2 FILLER_13_503 ();
 sg13g2_decap_8 FILLER_13_516 ();
 sg13g2_fill_2 FILLER_13_523 ();
 sg13g2_decap_4 FILLER_13_531 ();
 sg13g2_fill_1 FILLER_13_535 ();
 sg13g2_decap_4 FILLER_13_541 ();
 sg13g2_fill_2 FILLER_13_545 ();
 sg13g2_fill_2 FILLER_13_573 ();
 sg13g2_fill_1 FILLER_13_575 ();
 sg13g2_fill_2 FILLER_13_589 ();
 sg13g2_fill_1 FILLER_13_591 ();
 sg13g2_fill_1 FILLER_13_610 ();
 sg13g2_fill_2 FILLER_13_678 ();
 sg13g2_fill_1 FILLER_13_680 ();
 sg13g2_fill_2 FILLER_13_696 ();
 sg13g2_fill_1 FILLER_13_706 ();
 sg13g2_decap_4 FILLER_13_726 ();
 sg13g2_fill_1 FILLER_13_746 ();
 sg13g2_fill_2 FILLER_13_822 ();
 sg13g2_fill_2 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_4 FILLER_13_870 ();
 sg13g2_fill_2 FILLER_13_889 ();
 sg13g2_fill_1 FILLER_13_891 ();
 sg13g2_fill_2 FILLER_13_896 ();
 sg13g2_decap_8 FILLER_13_908 ();
 sg13g2_decap_8 FILLER_13_915 ();
 sg13g2_decap_8 FILLER_13_922 ();
 sg13g2_fill_1 FILLER_13_929 ();
 sg13g2_decap_8 FILLER_13_934 ();
 sg13g2_decap_4 FILLER_13_941 ();
 sg13g2_fill_1 FILLER_13_981 ();
 sg13g2_fill_1 FILLER_13_995 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_4 FILLER_13_1029 ();
 sg13g2_fill_1 FILLER_13_1033 ();
 sg13g2_decap_4 FILLER_13_1038 ();
 sg13g2_fill_2 FILLER_13_1042 ();
 sg13g2_decap_8 FILLER_13_1052 ();
 sg13g2_fill_2 FILLER_13_1059 ();
 sg13g2_fill_1 FILLER_13_1061 ();
 sg13g2_fill_2 FILLER_13_1070 ();
 sg13g2_decap_8 FILLER_13_1097 ();
 sg13g2_fill_1 FILLER_13_1104 ();
 sg13g2_decap_8 FILLER_13_1119 ();
 sg13g2_decap_8 FILLER_13_1126 ();
 sg13g2_decap_8 FILLER_13_1133 ();
 sg13g2_decap_8 FILLER_13_1140 ();
 sg13g2_decap_8 FILLER_13_1147 ();
 sg13g2_decap_8 FILLER_13_1154 ();
 sg13g2_decap_8 FILLER_13_1161 ();
 sg13g2_decap_8 FILLER_13_1168 ();
 sg13g2_decap_8 FILLER_13_1175 ();
 sg13g2_decap_8 FILLER_13_1182 ();
 sg13g2_decap_8 FILLER_13_1189 ();
 sg13g2_decap_8 FILLER_13_1196 ();
 sg13g2_decap_8 FILLER_13_1203 ();
 sg13g2_decap_8 FILLER_13_1210 ();
 sg13g2_decap_8 FILLER_13_1217 ();
 sg13g2_decap_8 FILLER_13_1224 ();
 sg13g2_decap_8 FILLER_13_1231 ();
 sg13g2_decap_8 FILLER_13_1238 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_decap_8 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_decap_8 FILLER_13_1280 ();
 sg13g2_decap_8 FILLER_13_1287 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1301 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_10 ();
 sg13g2_fill_2 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_20 ();
 sg13g2_fill_2 FILLER_14_24 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_decap_4 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_73 ();
 sg13g2_decap_8 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_decap_4 FILLER_14_148 ();
 sg13g2_decap_8 FILLER_14_156 ();
 sg13g2_decap_4 FILLER_14_163 ();
 sg13g2_fill_2 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_decap_4 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_250 ();
 sg13g2_decap_4 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_260 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_393 ();
 sg13g2_fill_2 FILLER_14_429 ();
 sg13g2_fill_1 FILLER_14_431 ();
 sg13g2_fill_1 FILLER_14_444 ();
 sg13g2_decap_8 FILLER_14_449 ();
 sg13g2_decap_4 FILLER_14_456 ();
 sg13g2_fill_2 FILLER_14_474 ();
 sg13g2_fill_1 FILLER_14_476 ();
 sg13g2_decap_4 FILLER_14_481 ();
 sg13g2_fill_1 FILLER_14_485 ();
 sg13g2_fill_2 FILLER_14_491 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_fill_1 FILLER_14_515 ();
 sg13g2_decap_8 FILLER_14_548 ();
 sg13g2_fill_2 FILLER_14_555 ();
 sg13g2_fill_1 FILLER_14_557 ();
 sg13g2_fill_2 FILLER_14_562 ();
 sg13g2_fill_1 FILLER_14_564 ();
 sg13g2_fill_2 FILLER_14_575 ();
 sg13g2_fill_1 FILLER_14_577 ();
 sg13g2_decap_4 FILLER_14_591 ();
 sg13g2_fill_2 FILLER_14_614 ();
 sg13g2_fill_1 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_635 ();
 sg13g2_decap_4 FILLER_14_673 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_decap_4 FILLER_14_716 ();
 sg13g2_fill_2 FILLER_14_731 ();
 sg13g2_fill_1 FILLER_14_733 ();
 sg13g2_decap_4 FILLER_14_751 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_fill_2 FILLER_14_767 ();
 sg13g2_fill_1 FILLER_14_769 ();
 sg13g2_decap_8 FILLER_14_778 ();
 sg13g2_fill_2 FILLER_14_785 ();
 sg13g2_fill_2 FILLER_14_791 ();
 sg13g2_fill_1 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_799 ();
 sg13g2_fill_2 FILLER_14_813 ();
 sg13g2_fill_1 FILLER_14_829 ();
 sg13g2_fill_1 FILLER_14_881 ();
 sg13g2_fill_1 FILLER_14_908 ();
 sg13g2_fill_2 FILLER_14_950 ();
 sg13g2_decap_4 FILLER_14_962 ();
 sg13g2_fill_1 FILLER_14_970 ();
 sg13g2_fill_2 FILLER_14_979 ();
 sg13g2_decap_8 FILLER_14_989 ();
 sg13g2_decap_4 FILLER_14_996 ();
 sg13g2_fill_2 FILLER_14_1000 ();
 sg13g2_fill_1 FILLER_14_1032 ();
 sg13g2_decap_8 FILLER_14_1120 ();
 sg13g2_decap_8 FILLER_14_1127 ();
 sg13g2_decap_8 FILLER_14_1134 ();
 sg13g2_decap_8 FILLER_14_1141 ();
 sg13g2_decap_8 FILLER_14_1148 ();
 sg13g2_decap_8 FILLER_14_1155 ();
 sg13g2_decap_8 FILLER_14_1162 ();
 sg13g2_decap_8 FILLER_14_1169 ();
 sg13g2_decap_8 FILLER_14_1176 ();
 sg13g2_decap_8 FILLER_14_1183 ();
 sg13g2_decap_8 FILLER_14_1190 ();
 sg13g2_decap_8 FILLER_14_1197 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_8 FILLER_14_1211 ();
 sg13g2_decap_8 FILLER_14_1218 ();
 sg13g2_decap_8 FILLER_14_1225 ();
 sg13g2_decap_8 FILLER_14_1232 ();
 sg13g2_decap_8 FILLER_14_1239 ();
 sg13g2_decap_8 FILLER_14_1246 ();
 sg13g2_decap_8 FILLER_14_1253 ();
 sg13g2_decap_8 FILLER_14_1260 ();
 sg13g2_decap_8 FILLER_14_1267 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_decap_4 FILLER_14_1309 ();
 sg13g2_fill_2 FILLER_14_1313 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_decap_4 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_decap_4 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_153 ();
 sg13g2_decap_4 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_decap_4 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_decap_4 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_decap_4 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_2 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_285 ();
 sg13g2_decap_4 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_15_350 ();
 sg13g2_fill_1 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_363 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_fill_2 FILLER_15_398 ();
 sg13g2_fill_1 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_419 ();
 sg13g2_fill_1 FILLER_15_447 ();
 sg13g2_fill_2 FILLER_15_464 ();
 sg13g2_fill_1 FILLER_15_466 ();
 sg13g2_decap_4 FILLER_15_494 ();
 sg13g2_decap_4 FILLER_15_532 ();
 sg13g2_fill_1 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_547 ();
 sg13g2_fill_2 FILLER_15_554 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_4 FILLER_15_571 ();
 sg13g2_fill_2 FILLER_15_587 ();
 sg13g2_fill_1 FILLER_15_589 ();
 sg13g2_decap_4 FILLER_15_598 ();
 sg13g2_fill_2 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_fill_2 FILLER_15_651 ();
 sg13g2_fill_1 FILLER_15_667 ();
 sg13g2_fill_1 FILLER_15_677 ();
 sg13g2_fill_1 FILLER_15_683 ();
 sg13g2_fill_2 FILLER_15_746 ();
 sg13g2_fill_1 FILLER_15_748 ();
 sg13g2_fill_2 FILLER_15_785 ();
 sg13g2_fill_1 FILLER_15_787 ();
 sg13g2_decap_4 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_fill_2 FILLER_15_866 ();
 sg13g2_fill_1 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_fill_2 FILLER_15_879 ();
 sg13g2_fill_1 FILLER_15_938 ();
 sg13g2_fill_2 FILLER_15_949 ();
 sg13g2_fill_1 FILLER_15_951 ();
 sg13g2_decap_8 FILLER_15_1003 ();
 sg13g2_fill_2 FILLER_15_1031 ();
 sg13g2_fill_1 FILLER_15_1033 ();
 sg13g2_decap_4 FILLER_15_1055 ();
 sg13g2_decap_4 FILLER_15_1074 ();
 sg13g2_fill_2 FILLER_15_1078 ();
 sg13g2_fill_2 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1093 ();
 sg13g2_decap_4 FILLER_15_1100 ();
 sg13g2_fill_1 FILLER_15_1104 ();
 sg13g2_decap_8 FILLER_15_1109 ();
 sg13g2_decap_8 FILLER_15_1116 ();
 sg13g2_decap_8 FILLER_15_1123 ();
 sg13g2_decap_8 FILLER_15_1130 ();
 sg13g2_decap_8 FILLER_15_1137 ();
 sg13g2_decap_8 FILLER_15_1144 ();
 sg13g2_decap_8 FILLER_15_1151 ();
 sg13g2_decap_8 FILLER_15_1158 ();
 sg13g2_decap_8 FILLER_15_1165 ();
 sg13g2_decap_8 FILLER_15_1172 ();
 sg13g2_decap_8 FILLER_15_1179 ();
 sg13g2_decap_8 FILLER_15_1186 ();
 sg13g2_decap_8 FILLER_15_1193 ();
 sg13g2_decap_8 FILLER_15_1200 ();
 sg13g2_decap_8 FILLER_15_1207 ();
 sg13g2_decap_8 FILLER_15_1214 ();
 sg13g2_decap_8 FILLER_15_1221 ();
 sg13g2_decap_8 FILLER_15_1228 ();
 sg13g2_decap_8 FILLER_15_1235 ();
 sg13g2_decap_8 FILLER_15_1242 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_decap_8 FILLER_15_1270 ();
 sg13g2_decap_8 FILLER_15_1277 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_fill_2 FILLER_15_1312 ();
 sg13g2_fill_1 FILLER_15_1314 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_10 ();
 sg13g2_fill_1 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_19 ();
 sg13g2_decap_8 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_decap_4 FILLER_16_66 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_252 ();
 sg13g2_fill_1 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_fill_2 FILLER_16_430 ();
 sg13g2_fill_2 FILLER_16_436 ();
 sg13g2_fill_1 FILLER_16_438 ();
 sg13g2_fill_2 FILLER_16_457 ();
 sg13g2_fill_1 FILLER_16_459 ();
 sg13g2_fill_1 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_498 ();
 sg13g2_fill_1 FILLER_16_505 ();
 sg13g2_fill_2 FILLER_16_511 ();
 sg13g2_fill_1 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_4 FILLER_16_525 ();
 sg13g2_fill_2 FILLER_16_565 ();
 sg13g2_fill_2 FILLER_16_588 ();
 sg13g2_fill_2 FILLER_16_606 ();
 sg13g2_fill_2 FILLER_16_615 ();
 sg13g2_fill_2 FILLER_16_661 ();
 sg13g2_fill_1 FILLER_16_671 ();
 sg13g2_fill_2 FILLER_16_692 ();
 sg13g2_decap_4 FILLER_16_726 ();
 sg13g2_decap_8 FILLER_16_755 ();
 sg13g2_decap_8 FILLER_16_762 ();
 sg13g2_decap_4 FILLER_16_769 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_4 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_813 ();
 sg13g2_fill_2 FILLER_16_820 ();
 sg13g2_fill_1 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_4 FILLER_16_877 ();
 sg13g2_fill_2 FILLER_16_881 ();
 sg13g2_decap_8 FILLER_16_909 ();
 sg13g2_decap_4 FILLER_16_916 ();
 sg13g2_fill_2 FILLER_16_920 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_fill_2 FILLER_16_944 ();
 sg13g2_fill_1 FILLER_16_961 ();
 sg13g2_decap_4 FILLER_16_966 ();
 sg13g2_fill_1 FILLER_16_970 ();
 sg13g2_decap_8 FILLER_16_1025 ();
 sg13g2_fill_2 FILLER_16_1032 ();
 sg13g2_decap_4 FILLER_16_1042 ();
 sg13g2_fill_1 FILLER_16_1046 ();
 sg13g2_decap_8 FILLER_16_1055 ();
 sg13g2_decap_8 FILLER_16_1062 ();
 sg13g2_decap_4 FILLER_16_1069 ();
 sg13g2_decap_4 FILLER_16_1091 ();
 sg13g2_fill_2 FILLER_16_1095 ();
 sg13g2_fill_1 FILLER_16_1111 ();
 sg13g2_fill_2 FILLER_16_1122 ();
 sg13g2_decap_8 FILLER_16_1128 ();
 sg13g2_decap_8 FILLER_16_1135 ();
 sg13g2_decap_8 FILLER_16_1142 ();
 sg13g2_decap_8 FILLER_16_1149 ();
 sg13g2_decap_8 FILLER_16_1156 ();
 sg13g2_decap_8 FILLER_16_1163 ();
 sg13g2_decap_8 FILLER_16_1170 ();
 sg13g2_decap_8 FILLER_16_1177 ();
 sg13g2_decap_8 FILLER_16_1184 ();
 sg13g2_decap_8 FILLER_16_1191 ();
 sg13g2_decap_8 FILLER_16_1198 ();
 sg13g2_decap_8 FILLER_16_1205 ();
 sg13g2_decap_8 FILLER_16_1212 ();
 sg13g2_decap_8 FILLER_16_1219 ();
 sg13g2_decap_8 FILLER_16_1226 ();
 sg13g2_decap_8 FILLER_16_1233 ();
 sg13g2_decap_8 FILLER_16_1240 ();
 sg13g2_decap_8 FILLER_16_1247 ();
 sg13g2_decap_8 FILLER_16_1254 ();
 sg13g2_decap_8 FILLER_16_1261 ();
 sg13g2_decap_8 FILLER_16_1268 ();
 sg13g2_decap_8 FILLER_16_1275 ();
 sg13g2_decap_8 FILLER_16_1282 ();
 sg13g2_decap_8 FILLER_16_1289 ();
 sg13g2_decap_8 FILLER_16_1296 ();
 sg13g2_decap_8 FILLER_16_1303 ();
 sg13g2_decap_4 FILLER_16_1310 ();
 sg13g2_fill_1 FILLER_16_1314 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_39 ();
 sg13g2_fill_1 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_decap_8 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_90 ();
 sg13g2_decap_8 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_decap_8 FILLER_17_148 ();
 sg13g2_decap_4 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_243 ();
 sg13g2_decap_4 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_4 FILLER_17_295 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_decap_4 FILLER_17_376 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_411 ();
 sg13g2_fill_2 FILLER_17_418 ();
 sg13g2_fill_1 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_439 ();
 sg13g2_fill_1 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_454 ();
 sg13g2_decap_8 FILLER_17_461 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_decap_8 FILLER_17_474 ();
 sg13g2_decap_8 FILLER_17_481 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_2 FILLER_17_542 ();
 sg13g2_fill_2 FILLER_17_568 ();
 sg13g2_fill_1 FILLER_17_570 ();
 sg13g2_decap_4 FILLER_17_588 ();
 sg13g2_decap_4 FILLER_17_602 ();
 sg13g2_fill_2 FILLER_17_606 ();
 sg13g2_fill_2 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_621 ();
 sg13g2_decap_8 FILLER_17_628 ();
 sg13g2_fill_1 FILLER_17_635 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_decap_8 FILLER_17_647 ();
 sg13g2_decap_4 FILLER_17_654 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_fill_2 FILLER_17_676 ();
 sg13g2_decap_4 FILLER_17_682 ();
 sg13g2_fill_2 FILLER_17_686 ();
 sg13g2_decap_4 FILLER_17_693 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_fill_1 FILLER_17_710 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_fill_1 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_734 ();
 sg13g2_fill_2 FILLER_17_741 ();
 sg13g2_fill_1 FILLER_17_743 ();
 sg13g2_fill_2 FILLER_17_788 ();
 sg13g2_fill_1 FILLER_17_806 ();
 sg13g2_decap_8 FILLER_17_886 ();
 sg13g2_fill_1 FILLER_17_893 ();
 sg13g2_fill_1 FILLER_17_898 ();
 sg13g2_fill_1 FILLER_17_935 ();
 sg13g2_fill_2 FILLER_17_946 ();
 sg13g2_decap_8 FILLER_17_972 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_4 FILLER_17_1001 ();
 sg13g2_fill_1 FILLER_17_1009 ();
 sg13g2_decap_8 FILLER_17_1014 ();
 sg13g2_decap_4 FILLER_17_1021 ();
 sg13g2_fill_2 FILLER_17_1025 ();
 sg13g2_fill_1 FILLER_17_1053 ();
 sg13g2_decap_4 FILLER_17_1062 ();
 sg13g2_fill_2 FILLER_17_1085 ();
 sg13g2_fill_1 FILLER_17_1087 ();
 sg13g2_decap_8 FILLER_17_1140 ();
 sg13g2_decap_8 FILLER_17_1147 ();
 sg13g2_decap_8 FILLER_17_1154 ();
 sg13g2_decap_8 FILLER_17_1161 ();
 sg13g2_decap_8 FILLER_17_1168 ();
 sg13g2_decap_8 FILLER_17_1175 ();
 sg13g2_decap_8 FILLER_17_1182 ();
 sg13g2_decap_8 FILLER_17_1189 ();
 sg13g2_decap_8 FILLER_17_1196 ();
 sg13g2_decap_8 FILLER_17_1203 ();
 sg13g2_decap_8 FILLER_17_1210 ();
 sg13g2_decap_8 FILLER_17_1217 ();
 sg13g2_decap_8 FILLER_17_1224 ();
 sg13g2_decap_8 FILLER_17_1231 ();
 sg13g2_decap_8 FILLER_17_1238 ();
 sg13g2_decap_8 FILLER_17_1245 ();
 sg13g2_decap_8 FILLER_17_1252 ();
 sg13g2_decap_8 FILLER_17_1259 ();
 sg13g2_decap_8 FILLER_17_1266 ();
 sg13g2_decap_8 FILLER_17_1273 ();
 sg13g2_decap_8 FILLER_17_1280 ();
 sg13g2_decap_8 FILLER_17_1287 ();
 sg13g2_decap_8 FILLER_17_1294 ();
 sg13g2_decap_8 FILLER_17_1301 ();
 sg13g2_decap_8 FILLER_17_1308 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_36 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_4 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_decap_4 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_decap_4 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_decap_4 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_fill_1 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_432 ();
 sg13g2_fill_1 FILLER_18_441 ();
 sg13g2_fill_1 FILLER_18_448 ();
 sg13g2_fill_2 FILLER_18_499 ();
 sg13g2_fill_2 FILLER_18_509 ();
 sg13g2_fill_1 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_517 ();
 sg13g2_decap_4 FILLER_18_524 ();
 sg13g2_fill_1 FILLER_18_528 ();
 sg13g2_fill_1 FILLER_18_538 ();
 sg13g2_fill_2 FILLER_18_562 ();
 sg13g2_fill_2 FILLER_18_584 ();
 sg13g2_fill_1 FILLER_18_586 ();
 sg13g2_decap_4 FILLER_18_600 ();
 sg13g2_decap_4 FILLER_18_624 ();
 sg13g2_fill_1 FILLER_18_628 ();
 sg13g2_fill_1 FILLER_18_681 ();
 sg13g2_decap_4 FILLER_18_687 ();
 sg13g2_fill_1 FILLER_18_691 ();
 sg13g2_decap_4 FILLER_18_702 ();
 sg13g2_fill_2 FILLER_18_706 ();
 sg13g2_fill_2 FILLER_18_718 ();
 sg13g2_fill_1 FILLER_18_720 ();
 sg13g2_fill_1 FILLER_18_725 ();
 sg13g2_decap_4 FILLER_18_745 ();
 sg13g2_fill_1 FILLER_18_749 ();
 sg13g2_decap_4 FILLER_18_753 ();
 sg13g2_fill_1 FILLER_18_757 ();
 sg13g2_fill_2 FILLER_18_794 ();
 sg13g2_decap_4 FILLER_18_799 ();
 sg13g2_fill_1 FILLER_18_803 ();
 sg13g2_decap_4 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_fill_1 FILLER_18_843 ();
 sg13g2_decap_4 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_858 ();
 sg13g2_decap_4 FILLER_18_863 ();
 sg13g2_fill_1 FILLER_18_867 ();
 sg13g2_fill_2 FILLER_18_877 ();
 sg13g2_decap_4 FILLER_18_884 ();
 sg13g2_fill_1 FILLER_18_888 ();
 sg13g2_decap_8 FILLER_18_909 ();
 sg13g2_decap_4 FILLER_18_916 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_fill_2 FILLER_18_948 ();
 sg13g2_decap_4 FILLER_18_953 ();
 sg13g2_fill_1 FILLER_18_957 ();
 sg13g2_decap_8 FILLER_18_1030 ();
 sg13g2_fill_1 FILLER_18_1037 ();
 sg13g2_decap_8 FILLER_18_1042 ();
 sg13g2_decap_4 FILLER_18_1049 ();
 sg13g2_fill_2 FILLER_18_1053 ();
 sg13g2_decap_8 FILLER_18_1068 ();
 sg13g2_decap_4 FILLER_18_1085 ();
 sg13g2_fill_2 FILLER_18_1108 ();
 sg13g2_fill_1 FILLER_18_1110 ();
 sg13g2_decap_8 FILLER_18_1121 ();
 sg13g2_fill_1 FILLER_18_1128 ();
 sg13g2_decap_8 FILLER_18_1132 ();
 sg13g2_decap_8 FILLER_18_1139 ();
 sg13g2_decap_8 FILLER_18_1146 ();
 sg13g2_decap_8 FILLER_18_1153 ();
 sg13g2_decap_8 FILLER_18_1160 ();
 sg13g2_decap_8 FILLER_18_1167 ();
 sg13g2_decap_8 FILLER_18_1174 ();
 sg13g2_decap_8 FILLER_18_1181 ();
 sg13g2_decap_8 FILLER_18_1188 ();
 sg13g2_decap_8 FILLER_18_1195 ();
 sg13g2_decap_8 FILLER_18_1202 ();
 sg13g2_decap_8 FILLER_18_1209 ();
 sg13g2_decap_8 FILLER_18_1216 ();
 sg13g2_decap_8 FILLER_18_1223 ();
 sg13g2_decap_8 FILLER_18_1230 ();
 sg13g2_decap_8 FILLER_18_1237 ();
 sg13g2_decap_8 FILLER_18_1244 ();
 sg13g2_decap_8 FILLER_18_1251 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_8 FILLER_18_1265 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_8 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1286 ();
 sg13g2_decap_8 FILLER_18_1293 ();
 sg13g2_decap_8 FILLER_18_1300 ();
 sg13g2_decap_8 FILLER_18_1307 ();
 sg13g2_fill_1 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_19 ();
 sg13g2_decap_4 FILLER_19_26 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_decap_8 FILLER_19_65 ();
 sg13g2_decap_8 FILLER_19_72 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_2 FILLER_19_107 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_decap_4 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_4 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_411 ();
 sg13g2_decap_4 FILLER_19_416 ();
 sg13g2_fill_1 FILLER_19_420 ();
 sg13g2_decap_4 FILLER_19_433 ();
 sg13g2_fill_1 FILLER_19_437 ();
 sg13g2_fill_2 FILLER_19_447 ();
 sg13g2_decap_8 FILLER_19_460 ();
 sg13g2_fill_2 FILLER_19_467 ();
 sg13g2_fill_1 FILLER_19_469 ();
 sg13g2_decap_4 FILLER_19_478 ();
 sg13g2_fill_1 FILLER_19_482 ();
 sg13g2_fill_2 FILLER_19_490 ();
 sg13g2_fill_1 FILLER_19_492 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_decap_4 FILLER_19_535 ();
 sg13g2_fill_1 FILLER_19_543 ();
 sg13g2_fill_2 FILLER_19_565 ();
 sg13g2_fill_1 FILLER_19_567 ();
 sg13g2_fill_2 FILLER_19_584 ();
 sg13g2_fill_1 FILLER_19_586 ();
 sg13g2_fill_1 FILLER_19_603 ();
 sg13g2_decap_4 FILLER_19_612 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_decap_4 FILLER_19_632 ();
 sg13g2_fill_1 FILLER_19_636 ();
 sg13g2_decap_4 FILLER_19_673 ();
 sg13g2_fill_2 FILLER_19_677 ();
 sg13g2_fill_2 FILLER_19_705 ();
 sg13g2_fill_1 FILLER_19_707 ();
 sg13g2_fill_1 FILLER_19_729 ();
 sg13g2_decap_8 FILLER_19_771 ();
 sg13g2_fill_1 FILLER_19_778 ();
 sg13g2_decap_4 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_4 FILLER_19_809 ();
 sg13g2_fill_1 FILLER_19_813 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_fill_1 FILLER_19_847 ();
 sg13g2_fill_1 FILLER_19_882 ();
 sg13g2_fill_2 FILLER_19_893 ();
 sg13g2_fill_1 FILLER_19_895 ();
 sg13g2_fill_2 FILLER_19_899 ();
 sg13g2_fill_1 FILLER_19_901 ();
 sg13g2_decap_4 FILLER_19_946 ();
 sg13g2_decap_8 FILLER_19_960 ();
 sg13g2_fill_2 FILLER_19_971 ();
 sg13g2_decap_4 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1003 ();
 sg13g2_fill_1 FILLER_19_1010 ();
 sg13g2_decap_4 FILLER_19_1025 ();
 sg13g2_fill_2 FILLER_19_1029 ();
 sg13g2_fill_2 FILLER_19_1035 ();
 sg13g2_fill_1 FILLER_19_1037 ();
 sg13g2_decap_8 FILLER_19_1059 ();
 sg13g2_fill_2 FILLER_19_1066 ();
 sg13g2_fill_2 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1139 ();
 sg13g2_decap_8 FILLER_19_1146 ();
 sg13g2_decap_8 FILLER_19_1153 ();
 sg13g2_decap_8 FILLER_19_1160 ();
 sg13g2_decap_8 FILLER_19_1167 ();
 sg13g2_decap_8 FILLER_19_1174 ();
 sg13g2_decap_8 FILLER_19_1181 ();
 sg13g2_decap_8 FILLER_19_1188 ();
 sg13g2_decap_8 FILLER_19_1195 ();
 sg13g2_decap_8 FILLER_19_1202 ();
 sg13g2_decap_8 FILLER_19_1209 ();
 sg13g2_decap_8 FILLER_19_1216 ();
 sg13g2_decap_8 FILLER_19_1223 ();
 sg13g2_decap_8 FILLER_19_1230 ();
 sg13g2_decap_8 FILLER_19_1237 ();
 sg13g2_decap_8 FILLER_19_1244 ();
 sg13g2_decap_8 FILLER_19_1251 ();
 sg13g2_decap_8 FILLER_19_1258 ();
 sg13g2_decap_8 FILLER_19_1265 ();
 sg13g2_decap_8 FILLER_19_1272 ();
 sg13g2_decap_8 FILLER_19_1279 ();
 sg13g2_decap_8 FILLER_19_1286 ();
 sg13g2_decap_8 FILLER_19_1293 ();
 sg13g2_decap_8 FILLER_19_1300 ();
 sg13g2_decap_8 FILLER_19_1307 ();
 sg13g2_fill_1 FILLER_19_1314 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_4 FILLER_20_38 ();
 sg13g2_decap_8 FILLER_20_73 ();
 sg13g2_decap_4 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_decap_4 FILLER_20_127 ();
 sg13g2_fill_2 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_decap_4 FILLER_20_349 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_4 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_431 ();
 sg13g2_fill_2 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_464 ();
 sg13g2_fill_2 FILLER_20_471 ();
 sg13g2_decap_4 FILLER_20_494 ();
 sg13g2_fill_1 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_526 ();
 sg13g2_fill_2 FILLER_20_533 ();
 sg13g2_decap_8 FILLER_20_544 ();
 sg13g2_fill_1 FILLER_20_551 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_4 FILLER_20_586 ();
 sg13g2_fill_1 FILLER_20_594 ();
 sg13g2_decap_8 FILLER_20_605 ();
 sg13g2_fill_1 FILLER_20_617 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_fill_1 FILLER_20_662 ();
 sg13g2_fill_2 FILLER_20_689 ();
 sg13g2_fill_1 FILLER_20_691 ();
 sg13g2_fill_2 FILLER_20_701 ();
 sg13g2_fill_2 FILLER_20_707 ();
 sg13g2_fill_1 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_fill_2 FILLER_20_734 ();
 sg13g2_fill_1 FILLER_20_736 ();
 sg13g2_decap_4 FILLER_20_749 ();
 sg13g2_fill_1 FILLER_20_794 ();
 sg13g2_fill_1 FILLER_20_831 ();
 sg13g2_fill_2 FILLER_20_842 ();
 sg13g2_fill_1 FILLER_20_844 ();
 sg13g2_fill_1 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_916 ();
 sg13g2_fill_1 FILLER_20_923 ();
 sg13g2_fill_2 FILLER_20_928 ();
 sg13g2_fill_1 FILLER_20_930 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_fill_2 FILLER_20_942 ();
 sg13g2_fill_1 FILLER_20_944 ();
 sg13g2_decap_4 FILLER_20_950 ();
 sg13g2_fill_2 FILLER_20_988 ();
 sg13g2_decap_8 FILLER_20_1088 ();
 sg13g2_decap_8 FILLER_20_1105 ();
 sg13g2_fill_2 FILLER_20_1122 ();
 sg13g2_decap_8 FILLER_20_1128 ();
 sg13g2_decap_8 FILLER_20_1135 ();
 sg13g2_decap_8 FILLER_20_1142 ();
 sg13g2_decap_8 FILLER_20_1149 ();
 sg13g2_decap_8 FILLER_20_1156 ();
 sg13g2_decap_8 FILLER_20_1163 ();
 sg13g2_decap_8 FILLER_20_1170 ();
 sg13g2_decap_8 FILLER_20_1177 ();
 sg13g2_decap_8 FILLER_20_1184 ();
 sg13g2_decap_8 FILLER_20_1191 ();
 sg13g2_decap_8 FILLER_20_1198 ();
 sg13g2_decap_8 FILLER_20_1205 ();
 sg13g2_decap_8 FILLER_20_1212 ();
 sg13g2_decap_8 FILLER_20_1219 ();
 sg13g2_decap_8 FILLER_20_1226 ();
 sg13g2_decap_8 FILLER_20_1233 ();
 sg13g2_decap_8 FILLER_20_1240 ();
 sg13g2_decap_8 FILLER_20_1247 ();
 sg13g2_decap_8 FILLER_20_1254 ();
 sg13g2_decap_8 FILLER_20_1261 ();
 sg13g2_decap_8 FILLER_20_1268 ();
 sg13g2_decap_8 FILLER_20_1275 ();
 sg13g2_decap_8 FILLER_20_1282 ();
 sg13g2_decap_8 FILLER_20_1289 ();
 sg13g2_decap_8 FILLER_20_1296 ();
 sg13g2_decap_8 FILLER_20_1303 ();
 sg13g2_decap_4 FILLER_20_1310 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_12 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_fill_2 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_decap_8 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_21_415 ();
 sg13g2_fill_1 FILLER_21_417 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_1 FILLER_21_430 ();
 sg13g2_fill_1 FILLER_21_437 ();
 sg13g2_decap_8 FILLER_21_443 ();
 sg13g2_fill_2 FILLER_21_450 ();
 sg13g2_fill_1 FILLER_21_452 ();
 sg13g2_fill_2 FILLER_21_473 ();
 sg13g2_fill_2 FILLER_21_479 ();
 sg13g2_fill_1 FILLER_21_481 ();
 sg13g2_fill_2 FILLER_21_487 ();
 sg13g2_fill_2 FILLER_21_511 ();
 sg13g2_fill_1 FILLER_21_513 ();
 sg13g2_fill_2 FILLER_21_519 ();
 sg13g2_fill_1 FILLER_21_544 ();
 sg13g2_fill_2 FILLER_21_553 ();
 sg13g2_fill_1 FILLER_21_555 ();
 sg13g2_fill_2 FILLER_21_569 ();
 sg13g2_fill_1 FILLER_21_571 ();
 sg13g2_fill_1 FILLER_21_628 ();
 sg13g2_decap_4 FILLER_21_669 ();
 sg13g2_fill_1 FILLER_21_673 ();
 sg13g2_decap_4 FILLER_21_678 ();
 sg13g2_fill_1 FILLER_21_682 ();
 sg13g2_decap_4 FILLER_21_688 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_4 FILLER_21_756 ();
 sg13g2_fill_1 FILLER_21_760 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_4 FILLER_21_783 ();
 sg13g2_fill_2 FILLER_21_787 ();
 sg13g2_decap_4 FILLER_21_799 ();
 sg13g2_fill_2 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_809 ();
 sg13g2_fill_1 FILLER_21_828 ();
 sg13g2_decap_4 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_fill_2 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_860 ();
 sg13g2_decap_4 FILLER_21_867 ();
 sg13g2_fill_2 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_888 ();
 sg13g2_decap_4 FILLER_21_949 ();
 sg13g2_fill_2 FILLER_21_963 ();
 sg13g2_fill_1 FILLER_21_965 ();
 sg13g2_decap_8 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_999 ();
 sg13g2_decap_4 FILLER_21_1006 ();
 sg13g2_fill_2 FILLER_21_1014 ();
 sg13g2_decap_4 FILLER_21_1036 ();
 sg13g2_fill_1 FILLER_21_1040 ();
 sg13g2_decap_8 FILLER_21_1062 ();
 sg13g2_decap_4 FILLER_21_1069 ();
 sg13g2_decap_4 FILLER_21_1077 ();
 sg13g2_fill_2 FILLER_21_1107 ();
 sg13g2_fill_1 FILLER_21_1109 ();
 sg13g2_decap_8 FILLER_21_1141 ();
 sg13g2_decap_8 FILLER_21_1148 ();
 sg13g2_decap_8 FILLER_21_1155 ();
 sg13g2_decap_8 FILLER_21_1162 ();
 sg13g2_decap_8 FILLER_21_1169 ();
 sg13g2_decap_8 FILLER_21_1176 ();
 sg13g2_decap_8 FILLER_21_1183 ();
 sg13g2_decap_8 FILLER_21_1190 ();
 sg13g2_decap_8 FILLER_21_1197 ();
 sg13g2_decap_8 FILLER_21_1204 ();
 sg13g2_decap_8 FILLER_21_1211 ();
 sg13g2_decap_8 FILLER_21_1218 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1239 ();
 sg13g2_decap_8 FILLER_21_1246 ();
 sg13g2_decap_8 FILLER_21_1253 ();
 sg13g2_decap_8 FILLER_21_1260 ();
 sg13g2_decap_8 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1274 ();
 sg13g2_decap_8 FILLER_21_1281 ();
 sg13g2_decap_8 FILLER_21_1288 ();
 sg13g2_decap_8 FILLER_21_1295 ();
 sg13g2_decap_8 FILLER_21_1302 ();
 sg13g2_decap_4 FILLER_21_1309 ();
 sg13g2_fill_2 FILLER_21_1313 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_19 ();
 sg13g2_fill_1 FILLER_22_23 ();
 sg13g2_fill_1 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_decap_8 FILLER_22_78 ();
 sg13g2_decap_4 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_decap_8 FILLER_22_139 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_8 FILLER_22_153 ();
 sg13g2_decap_4 FILLER_22_164 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_4 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_decap_4 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_4 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_22_434 ();
 sg13g2_fill_2 FILLER_22_447 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_2 FILLER_22_487 ();
 sg13g2_fill_1 FILLER_22_489 ();
 sg13g2_decap_4 FILLER_22_500 ();
 sg13g2_fill_2 FILLER_22_504 ();
 sg13g2_fill_2 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_fill_2 FILLER_22_543 ();
 sg13g2_fill_1 FILLER_22_545 ();
 sg13g2_fill_1 FILLER_22_556 ();
 sg13g2_decap_8 FILLER_22_568 ();
 sg13g2_fill_2 FILLER_22_575 ();
 sg13g2_fill_1 FILLER_22_577 ();
 sg13g2_decap_8 FILLER_22_583 ();
 sg13g2_decap_4 FILLER_22_590 ();
 sg13g2_decap_4 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_616 ();
 sg13g2_fill_2 FILLER_22_627 ();
 sg13g2_fill_2 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_647 ();
 sg13g2_fill_1 FILLER_22_654 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_fill_2 FILLER_22_667 ();
 sg13g2_fill_1 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_674 ();
 sg13g2_decap_4 FILLER_22_681 ();
 sg13g2_decap_4 FILLER_22_700 ();
 sg13g2_fill_1 FILLER_22_704 ();
 sg13g2_decap_4 FILLER_22_713 ();
 sg13g2_fill_1 FILLER_22_717 ();
 sg13g2_fill_2 FILLER_22_728 ();
 sg13g2_fill_1 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_fill_1 FILLER_22_752 ();
 sg13g2_decap_4 FILLER_22_789 ();
 sg13g2_fill_2 FILLER_22_793 ();
 sg13g2_fill_1 FILLER_22_850 ();
 sg13g2_decap_8 FILLER_22_856 ();
 sg13g2_fill_1 FILLER_22_878 ();
 sg13g2_fill_1 FILLER_22_889 ();
 sg13g2_decap_4 FILLER_22_910 ();
 sg13g2_fill_1 FILLER_22_914 ();
 sg13g2_fill_2 FILLER_22_982 ();
 sg13g2_fill_2 FILLER_22_1025 ();
 sg13g2_fill_2 FILLER_22_1058 ();
 sg13g2_fill_1 FILLER_22_1060 ();
 sg13g2_fill_2 FILLER_22_1087 ();
 sg13g2_fill_1 FILLER_22_1089 ();
 sg13g2_decap_8 FILLER_22_1104 ();
 sg13g2_decap_8 FILLER_22_1111 ();
 sg13g2_decap_8 FILLER_22_1118 ();
 sg13g2_fill_1 FILLER_22_1125 ();
 sg13g2_fill_2 FILLER_22_1130 ();
 sg13g2_decap_8 FILLER_22_1135 ();
 sg13g2_decap_8 FILLER_22_1142 ();
 sg13g2_decap_8 FILLER_22_1149 ();
 sg13g2_decap_8 FILLER_22_1156 ();
 sg13g2_decap_8 FILLER_22_1163 ();
 sg13g2_decap_8 FILLER_22_1170 ();
 sg13g2_decap_8 FILLER_22_1177 ();
 sg13g2_decap_8 FILLER_22_1184 ();
 sg13g2_decap_8 FILLER_22_1191 ();
 sg13g2_decap_8 FILLER_22_1198 ();
 sg13g2_decap_8 FILLER_22_1205 ();
 sg13g2_decap_8 FILLER_22_1212 ();
 sg13g2_decap_8 FILLER_22_1219 ();
 sg13g2_decap_8 FILLER_22_1226 ();
 sg13g2_decap_8 FILLER_22_1233 ();
 sg13g2_decap_8 FILLER_22_1240 ();
 sg13g2_decap_8 FILLER_22_1247 ();
 sg13g2_decap_8 FILLER_22_1254 ();
 sg13g2_decap_8 FILLER_22_1261 ();
 sg13g2_decap_8 FILLER_22_1268 ();
 sg13g2_decap_8 FILLER_22_1275 ();
 sg13g2_decap_8 FILLER_22_1282 ();
 sg13g2_decap_8 FILLER_22_1289 ();
 sg13g2_decap_8 FILLER_22_1296 ();
 sg13g2_decap_8 FILLER_22_1303 ();
 sg13g2_decap_4 FILLER_22_1310 ();
 sg13g2_fill_1 FILLER_22_1314 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_411 ();
 sg13g2_decap_4 FILLER_23_427 ();
 sg13g2_fill_2 FILLER_23_431 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_fill_1 FILLER_23_454 ();
 sg13g2_decap_4 FILLER_23_470 ();
 sg13g2_fill_2 FILLER_23_474 ();
 sg13g2_fill_2 FILLER_23_493 ();
 sg13g2_fill_2 FILLER_23_510 ();
 sg13g2_decap_4 FILLER_23_539 ();
 sg13g2_fill_1 FILLER_23_543 ();
 sg13g2_fill_2 FILLER_23_549 ();
 sg13g2_decap_8 FILLER_23_559 ();
 sg13g2_fill_2 FILLER_23_586 ();
 sg13g2_fill_1 FILLER_23_588 ();
 sg13g2_fill_2 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_619 ();
 sg13g2_fill_1 FILLER_23_648 ();
 sg13g2_fill_1 FILLER_23_685 ();
 sg13g2_decap_4 FILLER_23_707 ();
 sg13g2_fill_2 FILLER_23_711 ();
 sg13g2_fill_1 FILLER_23_717 ();
 sg13g2_fill_2 FILLER_23_728 ();
 sg13g2_fill_1 FILLER_23_746 ();
 sg13g2_decap_4 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_4 FILLER_23_770 ();
 sg13g2_decap_4 FILLER_23_814 ();
 sg13g2_fill_1 FILLER_23_818 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_4 FILLER_23_843 ();
 sg13g2_decap_4 FILLER_23_855 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_871 ();
 sg13g2_fill_2 FILLER_23_877 ();
 sg13g2_fill_1 FILLER_23_915 ();
 sg13g2_decap_8 FILLER_23_920 ();
 sg13g2_fill_2 FILLER_23_927 ();
 sg13g2_fill_1 FILLER_23_929 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_4 FILLER_23_963 ();
 sg13g2_fill_2 FILLER_23_971 ();
 sg13g2_decap_8 FILLER_23_990 ();
 sg13g2_decap_8 FILLER_23_997 ();
 sg13g2_decap_8 FILLER_23_1004 ();
 sg13g2_decap_8 FILLER_23_1015 ();
 sg13g2_decap_8 FILLER_23_1022 ();
 sg13g2_fill_2 FILLER_23_1029 ();
 sg13g2_fill_2 FILLER_23_1035 ();
 sg13g2_fill_1 FILLER_23_1042 ();
 sg13g2_decap_8 FILLER_23_1047 ();
 sg13g2_fill_2 FILLER_23_1054 ();
 sg13g2_fill_2 FILLER_23_1074 ();
 sg13g2_decap_4 FILLER_23_1088 ();
 sg13g2_fill_2 FILLER_23_1092 ();
 sg13g2_decap_8 FILLER_23_1120 ();
 sg13g2_decap_4 FILLER_23_1127 ();
 sg13g2_decap_8 FILLER_23_1135 ();
 sg13g2_decap_8 FILLER_23_1142 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1156 ();
 sg13g2_decap_8 FILLER_23_1163 ();
 sg13g2_decap_8 FILLER_23_1170 ();
 sg13g2_decap_8 FILLER_23_1177 ();
 sg13g2_decap_8 FILLER_23_1184 ();
 sg13g2_decap_8 FILLER_23_1191 ();
 sg13g2_decap_8 FILLER_23_1198 ();
 sg13g2_decap_8 FILLER_23_1205 ();
 sg13g2_decap_8 FILLER_23_1212 ();
 sg13g2_decap_8 FILLER_23_1219 ();
 sg13g2_decap_8 FILLER_23_1226 ();
 sg13g2_decap_8 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1240 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1261 ();
 sg13g2_decap_8 FILLER_23_1268 ();
 sg13g2_decap_8 FILLER_23_1275 ();
 sg13g2_decap_8 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_decap_8 FILLER_23_1296 ();
 sg13g2_decap_8 FILLER_23_1303 ();
 sg13g2_decap_4 FILLER_23_1310 ();
 sg13g2_fill_1 FILLER_23_1314 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_decap_4 FILLER_24_20 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_2 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_166 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_decap_4 FILLER_24_256 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_324 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_decap_4 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_fill_2 FILLER_24_359 ();
 sg13g2_decap_4 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_2 FILLER_24_378 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_fill_1 FILLER_24_427 ();
 sg13g2_fill_2 FILLER_24_442 ();
 sg13g2_fill_1 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_455 ();
 sg13g2_decap_4 FILLER_24_467 ();
 sg13g2_fill_2 FILLER_24_471 ();
 sg13g2_decap_4 FILLER_24_483 ();
 sg13g2_fill_1 FILLER_24_487 ();
 sg13g2_fill_1 FILLER_24_498 ();
 sg13g2_fill_2 FILLER_24_502 ();
 sg13g2_decap_4 FILLER_24_509 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_2 FILLER_24_520 ();
 sg13g2_fill_1 FILLER_24_522 ();
 sg13g2_fill_1 FILLER_24_548 ();
 sg13g2_fill_2 FILLER_24_573 ();
 sg13g2_decap_4 FILLER_24_587 ();
 sg13g2_fill_2 FILLER_24_591 ();
 sg13g2_decap_8 FILLER_24_617 ();
 sg13g2_decap_8 FILLER_24_624 ();
 sg13g2_fill_2 FILLER_24_631 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_decap_4 FILLER_24_668 ();
 sg13g2_fill_1 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_decap_4 FILLER_24_684 ();
 sg13g2_fill_1 FILLER_24_701 ();
 sg13g2_decap_4 FILLER_24_728 ();
 sg13g2_fill_1 FILLER_24_732 ();
 sg13g2_fill_1 FILLER_24_778 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_fill_2 FILLER_24_796 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_decap_4 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_881 ();
 sg13g2_decap_8 FILLER_24_898 ();
 sg13g2_fill_2 FILLER_24_955 ();
 sg13g2_decap_4 FILLER_24_967 ();
 sg13g2_fill_2 FILLER_24_971 ();
 sg13g2_fill_2 FILLER_24_988 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1033 ();
 sg13g2_fill_2 FILLER_24_1039 ();
 sg13g2_fill_1 FILLER_24_1041 ();
 sg13g2_decap_4 FILLER_24_1058 ();
 sg13g2_decap_4 FILLER_24_1067 ();
 sg13g2_decap_4 FILLER_24_1096 ();
 sg13g2_fill_2 FILLER_24_1100 ();
 sg13g2_fill_1 FILLER_24_1109 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1153 ();
 sg13g2_decap_8 FILLER_24_1160 ();
 sg13g2_decap_8 FILLER_24_1167 ();
 sg13g2_decap_8 FILLER_24_1174 ();
 sg13g2_decap_8 FILLER_24_1181 ();
 sg13g2_decap_8 FILLER_24_1188 ();
 sg13g2_decap_8 FILLER_24_1195 ();
 sg13g2_decap_8 FILLER_24_1202 ();
 sg13g2_decap_8 FILLER_24_1209 ();
 sg13g2_decap_8 FILLER_24_1216 ();
 sg13g2_decap_8 FILLER_24_1223 ();
 sg13g2_decap_8 FILLER_24_1230 ();
 sg13g2_decap_8 FILLER_24_1237 ();
 sg13g2_decap_8 FILLER_24_1244 ();
 sg13g2_decap_8 FILLER_24_1251 ();
 sg13g2_decap_8 FILLER_24_1258 ();
 sg13g2_decap_8 FILLER_24_1265 ();
 sg13g2_decap_8 FILLER_24_1272 ();
 sg13g2_decap_8 FILLER_24_1279 ();
 sg13g2_decap_8 FILLER_24_1286 ();
 sg13g2_decap_8 FILLER_24_1293 ();
 sg13g2_decap_8 FILLER_24_1300 ();
 sg13g2_decap_8 FILLER_24_1307 ();
 sg13g2_fill_1 FILLER_24_1314 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_decap_4 FILLER_25_66 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_decap_4 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_decap_4 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_271 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_decap_4 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_430 ();
 sg13g2_fill_2 FILLER_25_436 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_fill_2 FILLER_25_446 ();
 sg13g2_fill_1 FILLER_25_448 ();
 sg13g2_fill_2 FILLER_25_460 ();
 sg13g2_fill_1 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_472 ();
 sg13g2_fill_2 FILLER_25_488 ();
 sg13g2_fill_2 FILLER_25_507 ();
 sg13g2_decap_4 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_538 ();
 sg13g2_fill_1 FILLER_25_545 ();
 sg13g2_fill_2 FILLER_25_574 ();
 sg13g2_fill_1 FILLER_25_585 ();
 sg13g2_fill_2 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_591 ();
 sg13g2_decap_8 FILLER_25_596 ();
 sg13g2_fill_2 FILLER_25_603 ();
 sg13g2_decap_4 FILLER_25_688 ();
 sg13g2_fill_2 FILLER_25_720 ();
 sg13g2_decap_8 FILLER_25_726 ();
 sg13g2_fill_2 FILLER_25_733 ();
 sg13g2_fill_2 FILLER_25_750 ();
 sg13g2_fill_1 FILLER_25_752 ();
 sg13g2_fill_2 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_843 ();
 sg13g2_fill_2 FILLER_25_858 ();
 sg13g2_fill_2 FILLER_25_870 ();
 sg13g2_fill_1 FILLER_25_872 ();
 sg13g2_fill_1 FILLER_25_899 ();
 sg13g2_fill_2 FILLER_25_905 ();
 sg13g2_fill_1 FILLER_25_907 ();
 sg13g2_fill_2 FILLER_25_918 ();
 sg13g2_decap_8 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_931 ();
 sg13g2_fill_2 FILLER_25_938 ();
 sg13g2_fill_1 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_972 ();
 sg13g2_fill_1 FILLER_25_979 ();
 sg13g2_decap_4 FILLER_25_990 ();
 sg13g2_fill_2 FILLER_25_994 ();
 sg13g2_decap_4 FILLER_25_1009 ();
 sg13g2_fill_2 FILLER_25_1013 ();
 sg13g2_fill_2 FILLER_25_1045 ();
 sg13g2_fill_2 FILLER_25_1055 ();
 sg13g2_fill_1 FILLER_25_1080 ();
 sg13g2_fill_1 FILLER_25_1085 ();
 sg13g2_decap_8 FILLER_25_1103 ();
 sg13g2_fill_1 FILLER_25_1110 ();
 sg13g2_decap_8 FILLER_25_1147 ();
 sg13g2_decap_8 FILLER_25_1154 ();
 sg13g2_decap_8 FILLER_25_1161 ();
 sg13g2_decap_8 FILLER_25_1168 ();
 sg13g2_decap_8 FILLER_25_1175 ();
 sg13g2_decap_8 FILLER_25_1182 ();
 sg13g2_decap_8 FILLER_25_1189 ();
 sg13g2_decap_8 FILLER_25_1196 ();
 sg13g2_decap_8 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1210 ();
 sg13g2_decap_8 FILLER_25_1217 ();
 sg13g2_decap_8 FILLER_25_1224 ();
 sg13g2_decap_8 FILLER_25_1231 ();
 sg13g2_decap_8 FILLER_25_1238 ();
 sg13g2_decap_8 FILLER_25_1245 ();
 sg13g2_decap_8 FILLER_25_1252 ();
 sg13g2_decap_8 FILLER_25_1259 ();
 sg13g2_decap_8 FILLER_25_1266 ();
 sg13g2_decap_8 FILLER_25_1273 ();
 sg13g2_decap_8 FILLER_25_1280 ();
 sg13g2_decap_8 FILLER_25_1287 ();
 sg13g2_decap_8 FILLER_25_1294 ();
 sg13g2_decap_8 FILLER_25_1301 ();
 sg13g2_decap_8 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_25 ();
 sg13g2_fill_2 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_decap_4 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_decap_4 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_decap_4 FILLER_26_402 ();
 sg13g2_fill_2 FILLER_26_430 ();
 sg13g2_fill_1 FILLER_26_449 ();
 sg13g2_fill_2 FILLER_26_468 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_fill_1 FILLER_26_476 ();
 sg13g2_fill_2 FILLER_26_481 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_fill_2 FILLER_26_524 ();
 sg13g2_fill_1 FILLER_26_526 ();
 sg13g2_fill_2 FILLER_26_565 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_fill_1 FILLER_26_585 ();
 sg13g2_fill_1 FILLER_26_605 ();
 sg13g2_fill_1 FILLER_26_616 ();
 sg13g2_fill_2 FILLER_26_627 ();
 sg13g2_fill_1 FILLER_26_629 ();
 sg13g2_fill_2 FILLER_26_647 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_fill_2 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_703 ();
 sg13g2_fill_1 FILLER_26_710 ();
 sg13g2_decap_8 FILLER_26_745 ();
 sg13g2_decap_4 FILLER_26_752 ();
 sg13g2_fill_2 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_800 ();
 sg13g2_fill_2 FILLER_26_807 ();
 sg13g2_decap_4 FILLER_26_835 ();
 sg13g2_decap_4 FILLER_26_865 ();
 sg13g2_fill_2 FILLER_26_869 ();
 sg13g2_fill_2 FILLER_26_876 ();
 sg13g2_decap_8 FILLER_26_892 ();
 sg13g2_decap_8 FILLER_26_899 ();
 sg13g2_fill_2 FILLER_26_906 ();
 sg13g2_fill_1 FILLER_26_908 ();
 sg13g2_decap_8 FILLER_26_943 ();
 sg13g2_fill_1 FILLER_26_964 ();
 sg13g2_fill_1 FILLER_26_992 ();
 sg13g2_decap_8 FILLER_26_1029 ();
 sg13g2_decap_4 FILLER_26_1036 ();
 sg13g2_fill_1 FILLER_26_1040 ();
 sg13g2_decap_8 FILLER_26_1046 ();
 sg13g2_fill_1 FILLER_26_1053 ();
 sg13g2_decap_4 FILLER_26_1059 ();
 sg13g2_fill_1 FILLER_26_1063 ();
 sg13g2_decap_4 FILLER_26_1069 ();
 sg13g2_decap_8 FILLER_26_1078 ();
 sg13g2_fill_2 FILLER_26_1104 ();
 sg13g2_decap_8 FILLER_26_1116 ();
 sg13g2_fill_2 FILLER_26_1123 ();
 sg13g2_fill_1 FILLER_26_1125 ();
 sg13g2_fill_2 FILLER_26_1130 ();
 sg13g2_decap_8 FILLER_26_1136 ();
 sg13g2_decap_8 FILLER_26_1143 ();
 sg13g2_decap_8 FILLER_26_1150 ();
 sg13g2_decap_8 FILLER_26_1157 ();
 sg13g2_decap_8 FILLER_26_1164 ();
 sg13g2_decap_8 FILLER_26_1171 ();
 sg13g2_decap_8 FILLER_26_1178 ();
 sg13g2_decap_8 FILLER_26_1185 ();
 sg13g2_decap_8 FILLER_26_1192 ();
 sg13g2_decap_8 FILLER_26_1199 ();
 sg13g2_decap_8 FILLER_26_1206 ();
 sg13g2_decap_8 FILLER_26_1213 ();
 sg13g2_decap_8 FILLER_26_1220 ();
 sg13g2_decap_8 FILLER_26_1227 ();
 sg13g2_decap_8 FILLER_26_1234 ();
 sg13g2_decap_8 FILLER_26_1241 ();
 sg13g2_decap_8 FILLER_26_1248 ();
 sg13g2_decap_8 FILLER_26_1255 ();
 sg13g2_decap_8 FILLER_26_1262 ();
 sg13g2_decap_8 FILLER_26_1269 ();
 sg13g2_decap_8 FILLER_26_1276 ();
 sg13g2_decap_8 FILLER_26_1283 ();
 sg13g2_decap_8 FILLER_26_1290 ();
 sg13g2_decap_8 FILLER_26_1297 ();
 sg13g2_decap_8 FILLER_26_1304 ();
 sg13g2_decap_4 FILLER_26_1311 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_decap_4 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_decap_4 FILLER_27_193 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_4 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_decap_4 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_2 FILLER_27_431 ();
 sg13g2_decap_4 FILLER_27_458 ();
 sg13g2_decap_4 FILLER_27_468 ();
 sg13g2_fill_1 FILLER_27_472 ();
 sg13g2_fill_2 FILLER_27_481 ();
 sg13g2_fill_2 FILLER_27_489 ();
 sg13g2_fill_1 FILLER_27_491 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_4 FILLER_27_526 ();
 sg13g2_fill_2 FILLER_27_539 ();
 sg13g2_fill_2 FILLER_27_551 ();
 sg13g2_fill_1 FILLER_27_553 ();
 sg13g2_fill_2 FILLER_27_571 ();
 sg13g2_fill_2 FILLER_27_579 ();
 sg13g2_fill_1 FILLER_27_581 ();
 sg13g2_fill_2 FILLER_27_591 ();
 sg13g2_fill_1 FILLER_27_593 ();
 sg13g2_decap_4 FILLER_27_600 ();
 sg13g2_fill_2 FILLER_27_604 ();
 sg13g2_decap_4 FILLER_27_621 ();
 sg13g2_fill_2 FILLER_27_633 ();
 sg13g2_fill_1 FILLER_27_635 ();
 sg13g2_decap_4 FILLER_27_640 ();
 sg13g2_fill_1 FILLER_27_644 ();
 sg13g2_fill_1 FILLER_27_654 ();
 sg13g2_fill_1 FILLER_27_658 ();
 sg13g2_decap_4 FILLER_27_685 ();
 sg13g2_decap_8 FILLER_27_698 ();
 sg13g2_fill_2 FILLER_27_705 ();
 sg13g2_fill_1 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_723 ();
 sg13g2_fill_1 FILLER_27_730 ();
 sg13g2_fill_2 FILLER_27_738 ();
 sg13g2_decap_4 FILLER_27_748 ();
 sg13g2_fill_2 FILLER_27_760 ();
 sg13g2_fill_2 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_4 FILLER_27_833 ();
 sg13g2_fill_1 FILLER_27_837 ();
 sg13g2_fill_2 FILLER_27_846 ();
 sg13g2_fill_2 FILLER_27_908 ();
 sg13g2_fill_1 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_916 ();
 sg13g2_decap_4 FILLER_27_923 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_fill_1 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1006 ();
 sg13g2_decap_4 FILLER_27_1017 ();
 sg13g2_decap_8 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1092 ();
 sg13g2_decap_8 FILLER_27_1146 ();
 sg13g2_decap_8 FILLER_27_1153 ();
 sg13g2_decap_8 FILLER_27_1160 ();
 sg13g2_decap_8 FILLER_27_1167 ();
 sg13g2_decap_8 FILLER_27_1174 ();
 sg13g2_decap_8 FILLER_27_1181 ();
 sg13g2_decap_8 FILLER_27_1188 ();
 sg13g2_decap_8 FILLER_27_1195 ();
 sg13g2_decap_8 FILLER_27_1202 ();
 sg13g2_decap_8 FILLER_27_1209 ();
 sg13g2_decap_8 FILLER_27_1216 ();
 sg13g2_decap_8 FILLER_27_1223 ();
 sg13g2_decap_8 FILLER_27_1230 ();
 sg13g2_decap_8 FILLER_27_1237 ();
 sg13g2_decap_8 FILLER_27_1244 ();
 sg13g2_decap_8 FILLER_27_1251 ();
 sg13g2_decap_8 FILLER_27_1258 ();
 sg13g2_decap_8 FILLER_27_1265 ();
 sg13g2_decap_8 FILLER_27_1272 ();
 sg13g2_decap_8 FILLER_27_1279 ();
 sg13g2_decap_8 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1300 ();
 sg13g2_decap_8 FILLER_27_1307 ();
 sg13g2_fill_1 FILLER_27_1314 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_55 ();
 sg13g2_decap_8 FILLER_28_62 ();
 sg13g2_decap_4 FILLER_28_69 ();
 sg13g2_decap_4 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_fill_2 FILLER_28_343 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_4 FILLER_28_423 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_2 FILLER_28_434 ();
 sg13g2_fill_2 FILLER_28_441 ();
 sg13g2_fill_1 FILLER_28_443 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_fill_2 FILLER_28_460 ();
 sg13g2_fill_1 FILLER_28_462 ();
 sg13g2_decap_4 FILLER_28_488 ();
 sg13g2_fill_1 FILLER_28_492 ();
 sg13g2_fill_2 FILLER_28_528 ();
 sg13g2_fill_2 FILLER_28_548 ();
 sg13g2_fill_1 FILLER_28_550 ();
 sg13g2_fill_2 FILLER_28_559 ();
 sg13g2_fill_1 FILLER_28_561 ();
 sg13g2_fill_2 FILLER_28_576 ();
 sg13g2_fill_1 FILLER_28_578 ();
 sg13g2_fill_1 FILLER_28_603 ();
 sg13g2_fill_2 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_631 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_4 FILLER_28_673 ();
 sg13g2_fill_2 FILLER_28_677 ();
 sg13g2_decap_4 FILLER_28_698 ();
 sg13g2_fill_1 FILLER_28_746 ();
 sg13g2_decap_4 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_fill_2 FILLER_28_824 ();
 sg13g2_fill_1 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_fill_2 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_882 ();
 sg13g2_fill_2 FILLER_28_910 ();
 sg13g2_decap_4 FILLER_28_922 ();
 sg13g2_decap_4 FILLER_28_930 ();
 sg13g2_fill_1 FILLER_28_934 ();
 sg13g2_fill_2 FILLER_28_940 ();
 sg13g2_fill_1 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_952 ();
 sg13g2_decap_8 FILLER_28_959 ();
 sg13g2_decap_4 FILLER_28_966 ();
 sg13g2_fill_1 FILLER_28_970 ();
 sg13g2_fill_2 FILLER_28_979 ();
 sg13g2_fill_1 FILLER_28_981 ();
 sg13g2_fill_2 FILLER_28_1018 ();
 sg13g2_decap_8 FILLER_28_1041 ();
 sg13g2_fill_1 FILLER_28_1048 ();
 sg13g2_decap_4 FILLER_28_1061 ();
 sg13g2_decap_4 FILLER_28_1089 ();
 sg13g2_fill_2 FILLER_28_1111 ();
 sg13g2_fill_1 FILLER_28_1113 ();
 sg13g2_decap_8 FILLER_28_1154 ();
 sg13g2_decap_8 FILLER_28_1161 ();
 sg13g2_decap_8 FILLER_28_1168 ();
 sg13g2_decap_8 FILLER_28_1175 ();
 sg13g2_decap_8 FILLER_28_1182 ();
 sg13g2_decap_8 FILLER_28_1189 ();
 sg13g2_decap_8 FILLER_28_1196 ();
 sg13g2_decap_8 FILLER_28_1203 ();
 sg13g2_decap_8 FILLER_28_1210 ();
 sg13g2_decap_8 FILLER_28_1217 ();
 sg13g2_decap_8 FILLER_28_1224 ();
 sg13g2_decap_8 FILLER_28_1231 ();
 sg13g2_decap_8 FILLER_28_1238 ();
 sg13g2_decap_8 FILLER_28_1245 ();
 sg13g2_decap_8 FILLER_28_1252 ();
 sg13g2_decap_8 FILLER_28_1259 ();
 sg13g2_decap_8 FILLER_28_1266 ();
 sg13g2_decap_8 FILLER_28_1273 ();
 sg13g2_decap_8 FILLER_28_1280 ();
 sg13g2_decap_8 FILLER_28_1287 ();
 sg13g2_decap_8 FILLER_28_1294 ();
 sg13g2_decap_8 FILLER_28_1301 ();
 sg13g2_decap_8 FILLER_28_1308 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_25 ();
 sg13g2_fill_2 FILLER_29_29 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_92 ();
 sg13g2_decap_8 FILLER_29_99 ();
 sg13g2_decap_8 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_4 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_318 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_fill_1 FILLER_29_409 ();
 sg13g2_fill_1 FILLER_29_418 ();
 sg13g2_decap_4 FILLER_29_454 ();
 sg13g2_decap_4 FILLER_29_463 ();
 sg13g2_fill_2 FILLER_29_471 ();
 sg13g2_fill_1 FILLER_29_473 ();
 sg13g2_decap_4 FILLER_29_487 ();
 sg13g2_fill_1 FILLER_29_491 ();
 sg13g2_fill_2 FILLER_29_507 ();
 sg13g2_fill_2 FILLER_29_518 ();
 sg13g2_fill_2 FILLER_29_528 ();
 sg13g2_decap_8 FILLER_29_535 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_fill_1 FILLER_29_544 ();
 sg13g2_fill_2 FILLER_29_553 ();
 sg13g2_fill_2 FILLER_29_560 ();
 sg13g2_fill_1 FILLER_29_562 ();
 sg13g2_fill_2 FILLER_29_568 ();
 sg13g2_fill_1 FILLER_29_570 ();
 sg13g2_fill_2 FILLER_29_591 ();
 sg13g2_fill_1 FILLER_29_593 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_622 ();
 sg13g2_fill_1 FILLER_29_629 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_decap_4 FILLER_29_684 ();
 sg13g2_fill_2 FILLER_29_688 ();
 sg13g2_fill_1 FILLER_29_698 ();
 sg13g2_decap_8 FILLER_29_722 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_fill_1 FILLER_29_731 ();
 sg13g2_fill_2 FILLER_29_749 ();
 sg13g2_fill_1 FILLER_29_751 ();
 sg13g2_fill_2 FILLER_29_766 ();
 sg13g2_fill_1 FILLER_29_768 ();
 sg13g2_fill_2 FILLER_29_799 ();
 sg13g2_fill_1 FILLER_29_801 ();
 sg13g2_decap_8 FILLER_29_806 ();
 sg13g2_decap_8 FILLER_29_813 ();
 sg13g2_decap_4 FILLER_29_834 ();
 sg13g2_decap_4 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_866 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_fill_1 FILLER_29_914 ();
 sg13g2_fill_2 FILLER_29_946 ();
 sg13g2_fill_2 FILLER_29_992 ();
 sg13g2_fill_1 FILLER_29_994 ();
 sg13g2_decap_4 FILLER_29_1005 ();
 sg13g2_fill_1 FILLER_29_1009 ();
 sg13g2_decap_4 FILLER_29_1014 ();
 sg13g2_fill_2 FILLER_29_1018 ();
 sg13g2_decap_4 FILLER_29_1025 ();
 sg13g2_fill_2 FILLER_29_1029 ();
 sg13g2_fill_2 FILLER_29_1041 ();
 sg13g2_fill_1 FILLER_29_1043 ();
 sg13g2_fill_2 FILLER_29_1075 ();
 sg13g2_fill_2 FILLER_29_1082 ();
 sg13g2_fill_1 FILLER_29_1084 ();
 sg13g2_fill_1 FILLER_29_1111 ();
 sg13g2_fill_2 FILLER_29_1117 ();
 sg13g2_decap_8 FILLER_29_1145 ();
 sg13g2_decap_8 FILLER_29_1152 ();
 sg13g2_decap_8 FILLER_29_1159 ();
 sg13g2_decap_8 FILLER_29_1166 ();
 sg13g2_decap_8 FILLER_29_1173 ();
 sg13g2_decap_8 FILLER_29_1180 ();
 sg13g2_decap_8 FILLER_29_1187 ();
 sg13g2_decap_8 FILLER_29_1194 ();
 sg13g2_decap_8 FILLER_29_1201 ();
 sg13g2_decap_8 FILLER_29_1208 ();
 sg13g2_decap_8 FILLER_29_1215 ();
 sg13g2_decap_8 FILLER_29_1222 ();
 sg13g2_decap_8 FILLER_29_1229 ();
 sg13g2_decap_8 FILLER_29_1236 ();
 sg13g2_decap_8 FILLER_29_1243 ();
 sg13g2_decap_8 FILLER_29_1250 ();
 sg13g2_decap_8 FILLER_29_1257 ();
 sg13g2_decap_8 FILLER_29_1264 ();
 sg13g2_decap_8 FILLER_29_1271 ();
 sg13g2_decap_8 FILLER_29_1278 ();
 sg13g2_decap_8 FILLER_29_1285 ();
 sg13g2_decap_8 FILLER_29_1292 ();
 sg13g2_decap_8 FILLER_29_1299 ();
 sg13g2_decap_8 FILLER_29_1306 ();
 sg13g2_fill_2 FILLER_29_1313 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_16 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_decap_4 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_fill_1 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_decap_4 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_308 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_386 ();
 sg13g2_fill_2 FILLER_30_390 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_30_414 ();
 sg13g2_decap_8 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_453 ();
 sg13g2_decap_8 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_fill_1 FILLER_30_487 ();
 sg13g2_fill_2 FILLER_30_496 ();
 sg13g2_fill_1 FILLER_30_498 ();
 sg13g2_fill_2 FILLER_30_525 ();
 sg13g2_fill_1 FILLER_30_557 ();
 sg13g2_fill_2 FILLER_30_578 ();
 sg13g2_fill_1 FILLER_30_580 ();
 sg13g2_decap_8 FILLER_30_594 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_decap_8 FILLER_30_633 ();
 sg13g2_fill_1 FILLER_30_640 ();
 sg13g2_decap_8 FILLER_30_645 ();
 sg13g2_decap_4 FILLER_30_652 ();
 sg13g2_fill_2 FILLER_30_656 ();
 sg13g2_fill_1 FILLER_30_698 ();
 sg13g2_fill_2 FILLER_30_708 ();
 sg13g2_fill_1 FILLER_30_733 ();
 sg13g2_decap_8 FILLER_30_841 ();
 sg13g2_decap_4 FILLER_30_848 ();
 sg13g2_fill_1 FILLER_30_852 ();
 sg13g2_fill_2 FILLER_30_857 ();
 sg13g2_decap_4 FILLER_30_869 ();
 sg13g2_fill_1 FILLER_30_873 ();
 sg13g2_decap_4 FILLER_30_882 ();
 sg13g2_fill_2 FILLER_30_886 ();
 sg13g2_decap_4 FILLER_30_902 ();
 sg13g2_fill_1 FILLER_30_906 ();
 sg13g2_fill_2 FILLER_30_943 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_fill_1 FILLER_30_965 ();
 sg13g2_decap_4 FILLER_30_970 ();
 sg13g2_fill_1 FILLER_30_974 ();
 sg13g2_fill_2 FILLER_30_1042 ();
 sg13g2_fill_1 FILLER_30_1044 ();
 sg13g2_fill_2 FILLER_30_1054 ();
 sg13g2_fill_2 FILLER_30_1065 ();
 sg13g2_fill_1 FILLER_30_1082 ();
 sg13g2_fill_2 FILLER_30_1106 ();
 sg13g2_decap_8 FILLER_30_1139 ();
 sg13g2_decap_8 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1153 ();
 sg13g2_decap_8 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1167 ();
 sg13g2_decap_8 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_decap_8 FILLER_30_1188 ();
 sg13g2_decap_8 FILLER_30_1195 ();
 sg13g2_decap_8 FILLER_30_1202 ();
 sg13g2_decap_8 FILLER_30_1209 ();
 sg13g2_decap_8 FILLER_30_1216 ();
 sg13g2_decap_8 FILLER_30_1223 ();
 sg13g2_decap_8 FILLER_30_1230 ();
 sg13g2_decap_8 FILLER_30_1237 ();
 sg13g2_decap_8 FILLER_30_1244 ();
 sg13g2_decap_8 FILLER_30_1251 ();
 sg13g2_decap_8 FILLER_30_1258 ();
 sg13g2_decap_8 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1272 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_decap_8 FILLER_30_1286 ();
 sg13g2_decap_8 FILLER_30_1293 ();
 sg13g2_decap_8 FILLER_30_1300 ();
 sg13g2_decap_8 FILLER_30_1307 ();
 sg13g2_fill_1 FILLER_30_1314 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_decap_8 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_65 ();
 sg13g2_decap_4 FILLER_31_72 ();
 sg13g2_decap_4 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_decap_4 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_4 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_decap_4 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_439 ();
 sg13g2_fill_2 FILLER_31_453 ();
 sg13g2_fill_1 FILLER_31_485 ();
 sg13g2_decap_4 FILLER_31_507 ();
 sg13g2_fill_2 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_fill_1 FILLER_31_528 ();
 sg13g2_fill_2 FILLER_31_544 ();
 sg13g2_fill_1 FILLER_31_550 ();
 sg13g2_decap_8 FILLER_31_555 ();
 sg13g2_fill_2 FILLER_31_567 ();
 sg13g2_fill_1 FILLER_31_574 ();
 sg13g2_decap_4 FILLER_31_598 ();
 sg13g2_fill_2 FILLER_31_602 ();
 sg13g2_fill_1 FILLER_31_614 ();
 sg13g2_fill_2 FILLER_31_635 ();
 sg13g2_decap_4 FILLER_31_656 ();
 sg13g2_fill_2 FILLER_31_668 ();
 sg13g2_fill_1 FILLER_31_670 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_fill_1 FILLER_31_692 ();
 sg13g2_fill_1 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_fill_2 FILLER_31_775 ();
 sg13g2_fill_1 FILLER_31_777 ();
 sg13g2_decap_4 FILLER_31_788 ();
 sg13g2_fill_1 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_4 FILLER_31_808 ();
 sg13g2_fill_1 FILLER_31_812 ();
 sg13g2_fill_2 FILLER_31_828 ();
 sg13g2_decap_4 FILLER_31_838 ();
 sg13g2_decap_4 FILLER_31_868 ();
 sg13g2_fill_2 FILLER_31_872 ();
 sg13g2_decap_8 FILLER_31_918 ();
 sg13g2_fill_2 FILLER_31_925 ();
 sg13g2_fill_1 FILLER_31_927 ();
 sg13g2_decap_8 FILLER_31_932 ();
 sg13g2_fill_1 FILLER_31_939 ();
 sg13g2_fill_2 FILLER_31_954 ();
 sg13g2_fill_1 FILLER_31_956 ();
 sg13g2_decap_4 FILLER_31_975 ();
 sg13g2_fill_2 FILLER_31_979 ();
 sg13g2_fill_1 FILLER_31_993 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_8 FILLER_31_1009 ();
 sg13g2_decap_4 FILLER_31_1038 ();
 sg13g2_decap_8 FILLER_31_1059 ();
 sg13g2_fill_1 FILLER_31_1073 ();
 sg13g2_decap_4 FILLER_31_1094 ();
 sg13g2_decap_8 FILLER_31_1101 ();
 sg13g2_fill_1 FILLER_31_1108 ();
 sg13g2_fill_1 FILLER_31_1122 ();
 sg13g2_fill_2 FILLER_31_1127 ();
 sg13g2_fill_2 FILLER_31_1133 ();
 sg13g2_fill_1 FILLER_31_1135 ();
 sg13g2_decap_8 FILLER_31_1139 ();
 sg13g2_decap_8 FILLER_31_1146 ();
 sg13g2_decap_8 FILLER_31_1153 ();
 sg13g2_decap_8 FILLER_31_1160 ();
 sg13g2_decap_8 FILLER_31_1167 ();
 sg13g2_decap_8 FILLER_31_1174 ();
 sg13g2_decap_8 FILLER_31_1181 ();
 sg13g2_decap_8 FILLER_31_1188 ();
 sg13g2_decap_8 FILLER_31_1195 ();
 sg13g2_decap_8 FILLER_31_1202 ();
 sg13g2_decap_8 FILLER_31_1209 ();
 sg13g2_decap_8 FILLER_31_1216 ();
 sg13g2_decap_8 FILLER_31_1223 ();
 sg13g2_decap_8 FILLER_31_1230 ();
 sg13g2_decap_8 FILLER_31_1237 ();
 sg13g2_decap_8 FILLER_31_1244 ();
 sg13g2_decap_8 FILLER_31_1251 ();
 sg13g2_decap_8 FILLER_31_1258 ();
 sg13g2_decap_8 FILLER_31_1265 ();
 sg13g2_decap_8 FILLER_31_1272 ();
 sg13g2_decap_8 FILLER_31_1279 ();
 sg13g2_decap_8 FILLER_31_1286 ();
 sg13g2_decap_8 FILLER_31_1293 ();
 sg13g2_decap_8 FILLER_31_1300 ();
 sg13g2_decap_8 FILLER_31_1307 ();
 sg13g2_fill_1 FILLER_31_1314 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_1 FILLER_32_45 ();
 sg13g2_decap_4 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_145 ();
 sg13g2_decap_4 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_159 ();
 sg13g2_fill_2 FILLER_32_169 ();
 sg13g2_fill_1 FILLER_32_171 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_399 ();
 sg13g2_fill_1 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_415 ();
 sg13g2_fill_2 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_fill_1 FILLER_32_447 ();
 sg13g2_decap_4 FILLER_32_463 ();
 sg13g2_decap_8 FILLER_32_481 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_fill_2 FILLER_32_495 ();
 sg13g2_decap_8 FILLER_32_538 ();
 sg13g2_fill_2 FILLER_32_545 ();
 sg13g2_fill_1 FILLER_32_547 ();
 sg13g2_fill_2 FILLER_32_552 ();
 sg13g2_fill_2 FILLER_32_567 ();
 sg13g2_fill_1 FILLER_32_569 ();
 sg13g2_fill_2 FILLER_32_599 ();
 sg13g2_fill_1 FILLER_32_601 ();
 sg13g2_decap_4 FILLER_32_614 ();
 sg13g2_fill_1 FILLER_32_618 ();
 sg13g2_decap_4 FILLER_32_634 ();
 sg13g2_fill_1 FILLER_32_638 ();
 sg13g2_fill_2 FILLER_32_648 ();
 sg13g2_fill_1 FILLER_32_650 ();
 sg13g2_decap_4 FILLER_32_656 ();
 sg13g2_fill_2 FILLER_32_660 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_fill_2 FILLER_32_696 ();
 sg13g2_decap_4 FILLER_32_701 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_decap_4 FILLER_32_733 ();
 sg13g2_fill_1 FILLER_32_745 ();
 sg13g2_fill_1 FILLER_32_750 ();
 sg13g2_fill_2 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_761 ();
 sg13g2_fill_2 FILLER_32_780 ();
 sg13g2_fill_1 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_fill_2 FILLER_32_858 ();
 sg13g2_decap_4 FILLER_32_879 ();
 sg13g2_fill_1 FILLER_32_883 ();
 sg13g2_fill_1 FILLER_32_893 ();
 sg13g2_decap_4 FILLER_32_898 ();
 sg13g2_fill_2 FILLER_32_902 ();
 sg13g2_fill_1 FILLER_32_912 ();
 sg13g2_decap_8 FILLER_32_949 ();
 sg13g2_decap_8 FILLER_32_961 ();
 sg13g2_decap_4 FILLER_32_989 ();
 sg13g2_fill_2 FILLER_32_1029 ();
 sg13g2_fill_2 FILLER_32_1044 ();
 sg13g2_decap_4 FILLER_32_1072 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_8 FILLER_32_1169 ();
 sg13g2_decap_8 FILLER_32_1176 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1204 ();
 sg13g2_decap_8 FILLER_32_1211 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_decap_8 FILLER_32_1246 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_4 FILLER_32_1309 ();
 sg13g2_fill_2 FILLER_32_1313 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_23 ();
 sg13g2_decap_8 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_decap_4 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_decap_4 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_4 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_decap_4 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_414 ();
 sg13g2_decap_4 FILLER_33_423 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_decap_4 FILLER_33_439 ();
 sg13g2_fill_1 FILLER_33_443 ();
 sg13g2_fill_1 FILLER_33_449 ();
 sg13g2_decap_8 FILLER_33_454 ();
 sg13g2_decap_8 FILLER_33_461 ();
 sg13g2_fill_2 FILLER_33_468 ();
 sg13g2_fill_1 FILLER_33_470 ();
 sg13g2_fill_1 FILLER_33_481 ();
 sg13g2_decap_8 FILLER_33_494 ();
 sg13g2_decap_8 FILLER_33_501 ();
 sg13g2_fill_1 FILLER_33_508 ();
 sg13g2_decap_4 FILLER_33_519 ();
 sg13g2_fill_2 FILLER_33_523 ();
 sg13g2_fill_2 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_535 ();
 sg13g2_fill_2 FILLER_33_548 ();
 sg13g2_fill_1 FILLER_33_558 ();
 sg13g2_decap_4 FILLER_33_576 ();
 sg13g2_fill_1 FILLER_33_580 ();
 sg13g2_decap_8 FILLER_33_586 ();
 sg13g2_decap_4 FILLER_33_593 ();
 sg13g2_fill_1 FILLER_33_597 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_fill_1 FILLER_33_681 ();
 sg13g2_decap_4 FILLER_33_711 ();
 sg13g2_fill_1 FILLER_33_715 ();
 sg13g2_decap_8 FILLER_33_724 ();
 sg13g2_decap_4 FILLER_33_731 ();
 sg13g2_decap_4 FILLER_33_771 ();
 sg13g2_fill_2 FILLER_33_775 ();
 sg13g2_fill_2 FILLER_33_803 ();
 sg13g2_fill_2 FILLER_33_823 ();
 sg13g2_fill_1 FILLER_33_825 ();
 sg13g2_decap_4 FILLER_33_834 ();
 sg13g2_fill_1 FILLER_33_838 ();
 sg13g2_fill_2 FILLER_33_853 ();
 sg13g2_fill_1 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_fill_2 FILLER_33_868 ();
 sg13g2_fill_1 FILLER_33_870 ();
 sg13g2_decap_8 FILLER_33_881 ();
 sg13g2_decap_4 FILLER_33_888 ();
 sg13g2_fill_1 FILLER_33_892 ();
 sg13g2_fill_1 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_923 ();
 sg13g2_fill_1 FILLER_33_930 ();
 sg13g2_fill_1 FILLER_33_991 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_decap_8 FILLER_33_1007 ();
 sg13g2_fill_1 FILLER_33_1018 ();
 sg13g2_decap_8 FILLER_33_1062 ();
 sg13g2_fill_2 FILLER_33_1069 ();
 sg13g2_decap_8 FILLER_33_1096 ();
 sg13g2_fill_1 FILLER_33_1103 ();
 sg13g2_decap_4 FILLER_33_1107 ();
 sg13g2_decap_4 FILLER_33_1115 ();
 sg13g2_decap_8 FILLER_33_1123 ();
 sg13g2_decap_8 FILLER_33_1130 ();
 sg13g2_decap_8 FILLER_33_1137 ();
 sg13g2_decap_8 FILLER_33_1144 ();
 sg13g2_decap_8 FILLER_33_1151 ();
 sg13g2_decap_8 FILLER_33_1158 ();
 sg13g2_decap_8 FILLER_33_1165 ();
 sg13g2_decap_8 FILLER_33_1172 ();
 sg13g2_decap_8 FILLER_33_1179 ();
 sg13g2_decap_8 FILLER_33_1186 ();
 sg13g2_decap_8 FILLER_33_1193 ();
 sg13g2_decap_8 FILLER_33_1200 ();
 sg13g2_decap_8 FILLER_33_1207 ();
 sg13g2_decap_8 FILLER_33_1214 ();
 sg13g2_decap_8 FILLER_33_1221 ();
 sg13g2_decap_8 FILLER_33_1228 ();
 sg13g2_decap_8 FILLER_33_1235 ();
 sg13g2_decap_8 FILLER_33_1242 ();
 sg13g2_decap_8 FILLER_33_1249 ();
 sg13g2_decap_8 FILLER_33_1256 ();
 sg13g2_decap_8 FILLER_33_1263 ();
 sg13g2_decap_8 FILLER_33_1270 ();
 sg13g2_decap_8 FILLER_33_1277 ();
 sg13g2_decap_8 FILLER_33_1284 ();
 sg13g2_decap_8 FILLER_33_1291 ();
 sg13g2_decap_8 FILLER_33_1298 ();
 sg13g2_decap_8 FILLER_33_1305 ();
 sg13g2_fill_2 FILLER_33_1312 ();
 sg13g2_fill_1 FILLER_33_1314 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_101 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_132 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_222 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_decap_4 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_2 FILLER_34_444 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_4 FILLER_34_490 ();
 sg13g2_fill_1 FILLER_34_494 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_4 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_561 ();
 sg13g2_fill_2 FILLER_34_588 ();
 sg13g2_fill_1 FILLER_34_590 ();
 sg13g2_fill_2 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_598 ();
 sg13g2_fill_1 FILLER_34_603 ();
 sg13g2_fill_1 FILLER_34_609 ();
 sg13g2_decap_4 FILLER_34_619 ();
 sg13g2_fill_2 FILLER_34_623 ();
 sg13g2_fill_2 FILLER_34_629 ();
 sg13g2_fill_1 FILLER_34_631 ();
 sg13g2_fill_2 FILLER_34_646 ();
 sg13g2_fill_1 FILLER_34_648 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_fill_1 FILLER_34_665 ();
 sg13g2_decap_4 FILLER_34_671 ();
 sg13g2_fill_2 FILLER_34_680 ();
 sg13g2_fill_1 FILLER_34_694 ();
 sg13g2_fill_2 FILLER_34_720 ();
 sg13g2_fill_1 FILLER_34_722 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_fill_1 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_760 ();
 sg13g2_decap_8 FILLER_34_767 ();
 sg13g2_fill_2 FILLER_34_774 ();
 sg13g2_fill_2 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_fill_2 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_829 ();
 sg13g2_fill_1 FILLER_34_836 ();
 sg13g2_fill_2 FILLER_34_845 ();
 sg13g2_decap_4 FILLER_34_867 ();
 sg13g2_fill_2 FILLER_34_953 ();
 sg13g2_fill_1 FILLER_34_963 ();
 sg13g2_decap_8 FILLER_34_974 ();
 sg13g2_decap_4 FILLER_34_981 ();
 sg13g2_fill_1 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_1043 ();
 sg13g2_fill_2 FILLER_34_1050 ();
 sg13g2_fill_2 FILLER_34_1062 ();
 sg13g2_fill_1 FILLER_34_1064 ();
 sg13g2_fill_2 FILLER_34_1070 ();
 sg13g2_fill_2 FILLER_34_1087 ();
 sg13g2_decap_8 FILLER_34_1115 ();
 sg13g2_fill_2 FILLER_34_1122 ();
 sg13g2_decap_8 FILLER_34_1128 ();
 sg13g2_decap_8 FILLER_34_1135 ();
 sg13g2_decap_8 FILLER_34_1142 ();
 sg13g2_decap_8 FILLER_34_1149 ();
 sg13g2_decap_8 FILLER_34_1156 ();
 sg13g2_decap_8 FILLER_34_1163 ();
 sg13g2_decap_8 FILLER_34_1170 ();
 sg13g2_decap_8 FILLER_34_1177 ();
 sg13g2_decap_8 FILLER_34_1184 ();
 sg13g2_decap_8 FILLER_34_1191 ();
 sg13g2_decap_8 FILLER_34_1198 ();
 sg13g2_decap_8 FILLER_34_1205 ();
 sg13g2_decap_8 FILLER_34_1212 ();
 sg13g2_decap_8 FILLER_34_1219 ();
 sg13g2_decap_8 FILLER_34_1226 ();
 sg13g2_decap_8 FILLER_34_1233 ();
 sg13g2_decap_8 FILLER_34_1240 ();
 sg13g2_decap_8 FILLER_34_1247 ();
 sg13g2_decap_8 FILLER_34_1254 ();
 sg13g2_decap_8 FILLER_34_1261 ();
 sg13g2_decap_8 FILLER_34_1268 ();
 sg13g2_decap_8 FILLER_34_1275 ();
 sg13g2_decap_8 FILLER_34_1282 ();
 sg13g2_decap_8 FILLER_34_1289 ();
 sg13g2_decap_8 FILLER_34_1296 ();
 sg13g2_decap_8 FILLER_34_1303 ();
 sg13g2_decap_4 FILLER_34_1310 ();
 sg13g2_fill_1 FILLER_34_1314 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_decap_4 FILLER_35_22 ();
 sg13g2_decap_8 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_decap_4 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_35_334 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_decap_4 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_439 ();
 sg13g2_fill_1 FILLER_35_446 ();
 sg13g2_fill_1 FILLER_35_459 ();
 sg13g2_fill_2 FILLER_35_488 ();
 sg13g2_fill_1 FILLER_35_526 ();
 sg13g2_fill_2 FILLER_35_539 ();
 sg13g2_fill_2 FILLER_35_565 ();
 sg13g2_decap_4 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_583 ();
 sg13g2_fill_2 FILLER_35_609 ();
 sg13g2_fill_2 FILLER_35_615 ();
 sg13g2_fill_2 FILLER_35_639 ();
 sg13g2_fill_1 FILLER_35_671 ();
 sg13g2_fill_2 FILLER_35_696 ();
 sg13g2_fill_1 FILLER_35_703 ();
 sg13g2_fill_2 FILLER_35_709 ();
 sg13g2_fill_2 FILLER_35_721 ();
 sg13g2_fill_1 FILLER_35_723 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_fill_1 FILLER_35_736 ();
 sg13g2_fill_1 FILLER_35_781 ();
 sg13g2_decap_4 FILLER_35_829 ();
 sg13g2_fill_1 FILLER_35_841 ();
 sg13g2_fill_2 FILLER_35_892 ();
 sg13g2_fill_1 FILLER_35_894 ();
 sg13g2_decap_8 FILLER_35_904 ();
 sg13g2_decap_8 FILLER_35_911 ();
 sg13g2_decap_8 FILLER_35_922 ();
 sg13g2_decap_8 FILLER_35_929 ();
 sg13g2_decap_8 FILLER_35_1000 ();
 sg13g2_decap_8 FILLER_35_1011 ();
 sg13g2_decap_8 FILLER_35_1018 ();
 sg13g2_decap_8 FILLER_35_1025 ();
 sg13g2_decap_8 FILLER_35_1032 ();
 sg13g2_decap_4 FILLER_35_1039 ();
 sg13g2_fill_2 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1068 ();
 sg13g2_fill_1 FILLER_35_1070 ();
 sg13g2_decap_8 FILLER_35_1079 ();
 sg13g2_decap_8 FILLER_35_1086 ();
 sg13g2_decap_4 FILLER_35_1093 ();
 sg13g2_fill_2 FILLER_35_1111 ();
 sg13g2_decap_8 FILLER_35_1139 ();
 sg13g2_decap_8 FILLER_35_1146 ();
 sg13g2_decap_8 FILLER_35_1153 ();
 sg13g2_decap_8 FILLER_35_1160 ();
 sg13g2_decap_8 FILLER_35_1167 ();
 sg13g2_decap_8 FILLER_35_1174 ();
 sg13g2_decap_8 FILLER_35_1181 ();
 sg13g2_decap_8 FILLER_35_1188 ();
 sg13g2_decap_8 FILLER_35_1195 ();
 sg13g2_decap_8 FILLER_35_1202 ();
 sg13g2_decap_8 FILLER_35_1209 ();
 sg13g2_decap_8 FILLER_35_1216 ();
 sg13g2_decap_8 FILLER_35_1223 ();
 sg13g2_decap_8 FILLER_35_1230 ();
 sg13g2_decap_8 FILLER_35_1237 ();
 sg13g2_decap_8 FILLER_35_1244 ();
 sg13g2_decap_8 FILLER_35_1251 ();
 sg13g2_decap_8 FILLER_35_1258 ();
 sg13g2_decap_8 FILLER_35_1265 ();
 sg13g2_decap_8 FILLER_35_1272 ();
 sg13g2_decap_8 FILLER_35_1279 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_decap_8 FILLER_35_1293 ();
 sg13g2_decap_8 FILLER_35_1300 ();
 sg13g2_decap_8 FILLER_35_1307 ();
 sg13g2_fill_1 FILLER_35_1314 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_4 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_decap_4 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_282 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_4 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_423 ();
 sg13g2_decap_4 FILLER_36_432 ();
 sg13g2_fill_1 FILLER_36_448 ();
 sg13g2_decap_4 FILLER_36_460 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_decap_8 FILLER_36_474 ();
 sg13g2_fill_1 FILLER_36_481 ();
 sg13g2_fill_1 FILLER_36_496 ();
 sg13g2_fill_2 FILLER_36_504 ();
 sg13g2_fill_1 FILLER_36_506 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_fill_2 FILLER_36_532 ();
 sg13g2_decap_4 FILLER_36_551 ();
 sg13g2_fill_1 FILLER_36_555 ();
 sg13g2_fill_2 FILLER_36_568 ();
 sg13g2_fill_2 FILLER_36_583 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_decap_4 FILLER_36_591 ();
 sg13g2_fill_2 FILLER_36_595 ();
 sg13g2_decap_4 FILLER_36_602 ();
 sg13g2_fill_1 FILLER_36_606 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_fill_2 FILLER_36_643 ();
 sg13g2_fill_1 FILLER_36_645 ();
 sg13g2_fill_2 FILLER_36_651 ();
 sg13g2_decap_4 FILLER_36_657 ();
 sg13g2_decap_4 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_674 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_fill_2 FILLER_36_686 ();
 sg13g2_fill_1 FILLER_36_688 ();
 sg13g2_fill_1 FILLER_36_711 ();
 sg13g2_fill_2 FILLER_36_732 ();
 sg13g2_fill_2 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_744 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_decap_4 FILLER_36_764 ();
 sg13g2_fill_1 FILLER_36_768 ();
 sg13g2_fill_1 FILLER_36_787 ();
 sg13g2_fill_2 FILLER_36_802 ();
 sg13g2_fill_1 FILLER_36_804 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_fill_2 FILLER_36_816 ();
 sg13g2_fill_1 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_fill_1 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_fill_2 FILLER_36_890 ();
 sg13g2_fill_1 FILLER_36_892 ();
 sg13g2_fill_2 FILLER_36_903 ();
 sg13g2_decap_4 FILLER_36_915 ();
 sg13g2_fill_1 FILLER_36_919 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_fill_1 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_948 ();
 sg13g2_fill_2 FILLER_36_955 ();
 sg13g2_decap_8 FILLER_36_970 ();
 sg13g2_fill_2 FILLER_36_977 ();
 sg13g2_fill_2 FILLER_36_983 ();
 sg13g2_fill_2 FILLER_36_1016 ();
 sg13g2_fill_1 FILLER_36_1018 ();
 sg13g2_decap_8 FILLER_36_1034 ();
 sg13g2_fill_2 FILLER_36_1045 ();
 sg13g2_fill_1 FILLER_36_1047 ();
 sg13g2_decap_8 FILLER_36_1066 ();
 sg13g2_decap_8 FILLER_36_1073 ();
 sg13g2_decap_8 FILLER_36_1096 ();
 sg13g2_decap_8 FILLER_36_1103 ();
 sg13g2_fill_2 FILLER_36_1110 ();
 sg13g2_fill_1 FILLER_36_1112 ();
 sg13g2_decap_8 FILLER_36_1126 ();
 sg13g2_decap_8 FILLER_36_1133 ();
 sg13g2_decap_8 FILLER_36_1140 ();
 sg13g2_decap_8 FILLER_36_1147 ();
 sg13g2_decap_8 FILLER_36_1154 ();
 sg13g2_decap_8 FILLER_36_1161 ();
 sg13g2_decap_8 FILLER_36_1168 ();
 sg13g2_decap_8 FILLER_36_1175 ();
 sg13g2_decap_8 FILLER_36_1182 ();
 sg13g2_decap_8 FILLER_36_1189 ();
 sg13g2_decap_8 FILLER_36_1196 ();
 sg13g2_decap_8 FILLER_36_1203 ();
 sg13g2_decap_8 FILLER_36_1210 ();
 sg13g2_decap_8 FILLER_36_1217 ();
 sg13g2_decap_8 FILLER_36_1224 ();
 sg13g2_decap_8 FILLER_36_1231 ();
 sg13g2_decap_8 FILLER_36_1238 ();
 sg13g2_decap_8 FILLER_36_1245 ();
 sg13g2_decap_8 FILLER_36_1252 ();
 sg13g2_decap_8 FILLER_36_1259 ();
 sg13g2_decap_8 FILLER_36_1266 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_decap_8 FILLER_36_1280 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1294 ();
 sg13g2_decap_8 FILLER_36_1301 ();
 sg13g2_decap_8 FILLER_36_1308 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_18 ();
 sg13g2_decap_4 FILLER_37_22 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_75 ();
 sg13g2_fill_1 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_4 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_327 ();
 sg13g2_decap_4 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_decap_4 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_37_434 ();
 sg13g2_fill_2 FILLER_37_449 ();
 sg13g2_fill_2 FILLER_37_465 ();
 sg13g2_fill_1 FILLER_37_467 ();
 sg13g2_fill_2 FILLER_37_482 ();
 sg13g2_fill_1 FILLER_37_484 ();
 sg13g2_fill_2 FILLER_37_489 ();
 sg13g2_fill_1 FILLER_37_491 ();
 sg13g2_fill_2 FILLER_37_504 ();
 sg13g2_decap_4 FILLER_37_531 ();
 sg13g2_decap_4 FILLER_37_539 ();
 sg13g2_fill_1 FILLER_37_543 ();
 sg13g2_fill_2 FILLER_37_555 ();
 sg13g2_decap_4 FILLER_37_565 ();
 sg13g2_fill_2 FILLER_37_569 ();
 sg13g2_decap_8 FILLER_37_575 ();
 sg13g2_fill_1 FILLER_37_582 ();
 sg13g2_fill_1 FILLER_37_591 ();
 sg13g2_fill_2 FILLER_37_603 ();
 sg13g2_fill_1 FILLER_37_605 ();
 sg13g2_fill_2 FILLER_37_623 ();
 sg13g2_fill_1 FILLER_37_645 ();
 sg13g2_decap_4 FILLER_37_651 ();
 sg13g2_fill_2 FILLER_37_663 ();
 sg13g2_fill_1 FILLER_37_665 ();
 sg13g2_fill_1 FILLER_37_675 ();
 sg13g2_fill_2 FILLER_37_696 ();
 sg13g2_fill_1 FILLER_37_698 ();
 sg13g2_fill_1 FILLER_37_704 ();
 sg13g2_decap_4 FILLER_37_734 ();
 sg13g2_fill_2 FILLER_37_746 ();
 sg13g2_fill_1 FILLER_37_748 ();
 sg13g2_decap_4 FILLER_37_775 ();
 sg13g2_fill_2 FILLER_37_779 ();
 sg13g2_fill_2 FILLER_37_820 ();
 sg13g2_decap_8 FILLER_37_936 ();
 sg13g2_decap_8 FILLER_37_955 ();
 sg13g2_fill_2 FILLER_37_998 ();
 sg13g2_fill_1 FILLER_37_1000 ();
 sg13g2_fill_2 FILLER_37_1005 ();
 sg13g2_decap_8 FILLER_37_1059 ();
 sg13g2_fill_2 FILLER_37_1066 ();
 sg13g2_fill_2 FILLER_37_1084 ();
 sg13g2_decap_8 FILLER_37_1129 ();
 sg13g2_decap_8 FILLER_37_1136 ();
 sg13g2_decap_8 FILLER_37_1143 ();
 sg13g2_decap_8 FILLER_37_1150 ();
 sg13g2_decap_8 FILLER_37_1157 ();
 sg13g2_decap_8 FILLER_37_1164 ();
 sg13g2_decap_8 FILLER_37_1171 ();
 sg13g2_decap_8 FILLER_37_1178 ();
 sg13g2_decap_8 FILLER_37_1185 ();
 sg13g2_decap_8 FILLER_37_1192 ();
 sg13g2_decap_8 FILLER_37_1199 ();
 sg13g2_decap_8 FILLER_37_1206 ();
 sg13g2_decap_8 FILLER_37_1213 ();
 sg13g2_decap_8 FILLER_37_1220 ();
 sg13g2_decap_8 FILLER_37_1227 ();
 sg13g2_decap_8 FILLER_37_1234 ();
 sg13g2_decap_8 FILLER_37_1241 ();
 sg13g2_decap_8 FILLER_37_1248 ();
 sg13g2_decap_8 FILLER_37_1255 ();
 sg13g2_decap_8 FILLER_37_1262 ();
 sg13g2_decap_8 FILLER_37_1269 ();
 sg13g2_decap_8 FILLER_37_1276 ();
 sg13g2_decap_8 FILLER_37_1283 ();
 sg13g2_decap_8 FILLER_37_1290 ();
 sg13g2_decap_8 FILLER_37_1297 ();
 sg13g2_decap_8 FILLER_37_1304 ();
 sg13g2_decap_4 FILLER_37_1311 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_1 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_235 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_288 ();
 sg13g2_decap_4 FILLER_38_313 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_decap_4 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_432 ();
 sg13g2_fill_2 FILLER_38_436 ();
 sg13g2_decap_4 FILLER_38_446 ();
 sg13g2_fill_1 FILLER_38_459 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_fill_2 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_495 ();
 sg13g2_decap_8 FILLER_38_502 ();
 sg13g2_fill_1 FILLER_38_509 ();
 sg13g2_fill_2 FILLER_38_523 ();
 sg13g2_fill_1 FILLER_38_555 ();
 sg13g2_decap_4 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_590 ();
 sg13g2_decap_4 FILLER_38_600 ();
 sg13g2_decap_4 FILLER_38_613 ();
 sg13g2_fill_1 FILLER_38_617 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_4 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_634 ();
 sg13g2_decap_4 FILLER_38_653 ();
 sg13g2_fill_2 FILLER_38_657 ();
 sg13g2_fill_1 FILLER_38_663 ();
 sg13g2_fill_2 FILLER_38_679 ();
 sg13g2_decap_4 FILLER_38_685 ();
 sg13g2_fill_1 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_713 ();
 sg13g2_fill_2 FILLER_38_720 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_decap_8 FILLER_38_744 ();
 sg13g2_fill_2 FILLER_38_780 ();
 sg13g2_decap_8 FILLER_38_790 ();
 sg13g2_decap_8 FILLER_38_797 ();
 sg13g2_decap_4 FILLER_38_804 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_fill_2 FILLER_38_830 ();
 sg13g2_fill_1 FILLER_38_832 ();
 sg13g2_fill_2 FILLER_38_841 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_4 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_871 ();
 sg13g2_fill_2 FILLER_38_878 ();
 sg13g2_fill_2 FILLER_38_885 ();
 sg13g2_fill_1 FILLER_38_887 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_fill_2 FILLER_38_903 ();
 sg13g2_fill_1 FILLER_38_905 ();
 sg13g2_decap_8 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_4 FILLER_38_928 ();
 sg13g2_fill_2 FILLER_38_932 ();
 sg13g2_fill_1 FILLER_38_942 ();
 sg13g2_decap_4 FILLER_38_977 ();
 sg13g2_fill_2 FILLER_38_981 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_fill_2 FILLER_38_1001 ();
 sg13g2_decap_4 FILLER_38_1013 ();
 sg13g2_fill_1 FILLER_38_1017 ();
 sg13g2_fill_1 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_38_1032 ();
 sg13g2_decap_4 FILLER_38_1070 ();
 sg13g2_fill_1 FILLER_38_1074 ();
 sg13g2_fill_2 FILLER_38_1111 ();
 sg13g2_decap_8 FILLER_38_1117 ();
 sg13g2_decap_8 FILLER_38_1124 ();
 sg13g2_decap_8 FILLER_38_1131 ();
 sg13g2_decap_8 FILLER_38_1138 ();
 sg13g2_decap_8 FILLER_38_1145 ();
 sg13g2_decap_8 FILLER_38_1152 ();
 sg13g2_decap_8 FILLER_38_1159 ();
 sg13g2_decap_8 FILLER_38_1166 ();
 sg13g2_decap_8 FILLER_38_1173 ();
 sg13g2_decap_8 FILLER_38_1180 ();
 sg13g2_decap_8 FILLER_38_1187 ();
 sg13g2_decap_8 FILLER_38_1194 ();
 sg13g2_decap_8 FILLER_38_1201 ();
 sg13g2_decap_8 FILLER_38_1208 ();
 sg13g2_decap_8 FILLER_38_1215 ();
 sg13g2_decap_8 FILLER_38_1222 ();
 sg13g2_decap_8 FILLER_38_1229 ();
 sg13g2_decap_8 FILLER_38_1236 ();
 sg13g2_decap_8 FILLER_38_1243 ();
 sg13g2_decap_8 FILLER_38_1250 ();
 sg13g2_decap_8 FILLER_38_1257 ();
 sg13g2_decap_8 FILLER_38_1264 ();
 sg13g2_decap_8 FILLER_38_1271 ();
 sg13g2_decap_8 FILLER_38_1278 ();
 sg13g2_decap_8 FILLER_38_1285 ();
 sg13g2_decap_8 FILLER_38_1292 ();
 sg13g2_decap_8 FILLER_38_1299 ();
 sg13g2_decap_8 FILLER_38_1306 ();
 sg13g2_fill_2 FILLER_38_1313 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_23 ();
 sg13g2_decap_8 FILLER_39_34 ();
 sg13g2_fill_2 FILLER_39_41 ();
 sg13g2_fill_1 FILLER_39_48 ();
 sg13g2_decap_8 FILLER_39_75 ();
 sg13g2_fill_1 FILLER_39_82 ();
 sg13g2_decap_8 FILLER_39_103 ();
 sg13g2_decap_4 FILLER_39_110 ();
 sg13g2_fill_2 FILLER_39_118 ();
 sg13g2_fill_1 FILLER_39_120 ();
 sg13g2_decap_8 FILLER_39_129 ();
 sg13g2_decap_4 FILLER_39_136 ();
 sg13g2_fill_2 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_150 ();
 sg13g2_fill_2 FILLER_39_177 ();
 sg13g2_decap_8 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_decap_4 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_248 ();
 sg13g2_fill_1 FILLER_39_250 ();
 sg13g2_decap_4 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_decap_4 FILLER_39_281 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_339 ();
 sg13g2_fill_2 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_397 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_fill_1 FILLER_39_456 ();
 sg13g2_fill_1 FILLER_39_471 ();
 sg13g2_decap_8 FILLER_39_481 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_fill_1 FILLER_39_505 ();
 sg13g2_fill_1 FILLER_39_522 ();
 sg13g2_fill_2 FILLER_39_528 ();
 sg13g2_fill_1 FILLER_39_530 ();
 sg13g2_fill_2 FILLER_39_535 ();
 sg13g2_fill_2 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_551 ();
 sg13g2_fill_2 FILLER_39_564 ();
 sg13g2_fill_1 FILLER_39_566 ();
 sg13g2_fill_2 FILLER_39_584 ();
 sg13g2_fill_1 FILLER_39_586 ();
 sg13g2_fill_2 FILLER_39_597 ();
 sg13g2_fill_2 FILLER_39_614 ();
 sg13g2_fill_1 FILLER_39_616 ();
 sg13g2_decap_4 FILLER_39_637 ();
 sg13g2_decap_4 FILLER_39_645 ();
 sg13g2_fill_2 FILLER_39_667 ();
 sg13g2_fill_2 FILLER_39_673 ();
 sg13g2_fill_1 FILLER_39_684 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_fill_2 FILLER_39_702 ();
 sg13g2_decap_4 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_734 ();
 sg13g2_decap_4 FILLER_39_754 ();
 sg13g2_fill_1 FILLER_39_758 ();
 sg13g2_decap_4 FILLER_39_790 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_fill_2 FILLER_39_831 ();
 sg13g2_fill_1 FILLER_39_833 ();
 sg13g2_fill_2 FILLER_39_838 ();
 sg13g2_fill_1 FILLER_39_840 ();
 sg13g2_fill_1 FILLER_39_850 ();
 sg13g2_fill_1 FILLER_39_860 ();
 sg13g2_decap_4 FILLER_39_865 ();
 sg13g2_decap_4 FILLER_39_956 ();
 sg13g2_fill_2 FILLER_39_973 ();
 sg13g2_fill_1 FILLER_39_975 ();
 sg13g2_decap_8 FILLER_39_981 ();
 sg13g2_decap_4 FILLER_39_988 ();
 sg13g2_fill_2 FILLER_39_992 ();
 sg13g2_decap_8 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1019 ();
 sg13g2_fill_1 FILLER_39_1026 ();
 sg13g2_decap_8 FILLER_39_1036 ();
 sg13g2_decap_8 FILLER_39_1043 ();
 sg13g2_fill_1 FILLER_39_1054 ();
 sg13g2_fill_1 FILLER_39_1065 ();
 sg13g2_decap_4 FILLER_39_1096 ();
 sg13g2_fill_2 FILLER_39_1100 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_decap_8 FILLER_39_1149 ();
 sg13g2_decap_8 FILLER_39_1156 ();
 sg13g2_decap_8 FILLER_39_1163 ();
 sg13g2_decap_8 FILLER_39_1170 ();
 sg13g2_decap_8 FILLER_39_1177 ();
 sg13g2_decap_8 FILLER_39_1184 ();
 sg13g2_decap_8 FILLER_39_1191 ();
 sg13g2_decap_8 FILLER_39_1198 ();
 sg13g2_decap_8 FILLER_39_1205 ();
 sg13g2_decap_8 FILLER_39_1212 ();
 sg13g2_decap_8 FILLER_39_1219 ();
 sg13g2_decap_8 FILLER_39_1226 ();
 sg13g2_decap_8 FILLER_39_1233 ();
 sg13g2_decap_8 FILLER_39_1240 ();
 sg13g2_decap_8 FILLER_39_1247 ();
 sg13g2_decap_8 FILLER_39_1254 ();
 sg13g2_decap_8 FILLER_39_1261 ();
 sg13g2_decap_8 FILLER_39_1268 ();
 sg13g2_decap_8 FILLER_39_1275 ();
 sg13g2_decap_8 FILLER_39_1282 ();
 sg13g2_decap_8 FILLER_39_1289 ();
 sg13g2_decap_8 FILLER_39_1296 ();
 sg13g2_decap_8 FILLER_39_1303 ();
 sg13g2_decap_4 FILLER_39_1310 ();
 sg13g2_fill_1 FILLER_39_1314 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_18 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_fill_1 FILLER_40_130 ();
 sg13g2_fill_1 FILLER_40_162 ();
 sg13g2_fill_2 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_267 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_decap_4 FILLER_40_279 ();
 sg13g2_decap_4 FILLER_40_295 ();
 sg13g2_fill_1 FILLER_40_299 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_decap_4 FILLER_40_317 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_346 ();
 sg13g2_decap_4 FILLER_40_379 ();
 sg13g2_fill_2 FILLER_40_383 ();
 sg13g2_decap_4 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_fill_2 FILLER_40_413 ();
 sg13g2_fill_1 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_424 ();
 sg13g2_decap_4 FILLER_40_431 ();
 sg13g2_fill_2 FILLER_40_444 ();
 sg13g2_fill_1 FILLER_40_446 ();
 sg13g2_fill_1 FILLER_40_485 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_fill_1 FILLER_40_531 ();
 sg13g2_decap_8 FILLER_40_552 ();
 sg13g2_fill_1 FILLER_40_559 ();
 sg13g2_decap_8 FILLER_40_565 ();
 sg13g2_decap_8 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_596 ();
 sg13g2_fill_2 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_612 ();
 sg13g2_decap_8 FILLER_40_619 ();
 sg13g2_fill_2 FILLER_40_630 ();
 sg13g2_fill_1 FILLER_40_632 ();
 sg13g2_decap_4 FILLER_40_650 ();
 sg13g2_fill_1 FILLER_40_654 ();
 sg13g2_fill_2 FILLER_40_660 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_fill_1 FILLER_40_682 ();
 sg13g2_decap_4 FILLER_40_688 ();
 sg13g2_fill_2 FILLER_40_706 ();
 sg13g2_decap_8 FILLER_40_732 ();
 sg13g2_decap_4 FILLER_40_739 ();
 sg13g2_fill_1 FILLER_40_743 ();
 sg13g2_decap_4 FILLER_40_757 ();
 sg13g2_fill_2 FILLER_40_761 ();
 sg13g2_decap_4 FILLER_40_775 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_fill_1 FILLER_40_786 ();
 sg13g2_fill_2 FILLER_40_821 ();
 sg13g2_fill_2 FILLER_40_849 ();
 sg13g2_decap_4 FILLER_40_877 ();
 sg13g2_fill_1 FILLER_40_881 ();
 sg13g2_decap_8 FILLER_40_891 ();
 sg13g2_decap_4 FILLER_40_898 ();
 sg13g2_fill_1 FILLER_40_906 ();
 sg13g2_decap_4 FILLER_40_919 ();
 sg13g2_fill_2 FILLER_40_923 ();
 sg13g2_fill_1 FILLER_40_934 ();
 sg13g2_fill_2 FILLER_40_1043 ();
 sg13g2_fill_1 FILLER_40_1045 ();
 sg13g2_decap_8 FILLER_40_1051 ();
 sg13g2_fill_1 FILLER_40_1058 ();
 sg13g2_decap_8 FILLER_40_1063 ();
 sg13g2_fill_2 FILLER_40_1070 ();
 sg13g2_fill_1 FILLER_40_1072 ();
 sg13g2_fill_2 FILLER_40_1085 ();
 sg13g2_fill_1 FILLER_40_1092 ();
 sg13g2_decap_4 FILLER_40_1101 ();
 sg13g2_fill_2 FILLER_40_1105 ();
 sg13g2_fill_1 FILLER_40_1112 ();
 sg13g2_decap_8 FILLER_40_1121 ();
 sg13g2_decap_8 FILLER_40_1128 ();
 sg13g2_decap_8 FILLER_40_1135 ();
 sg13g2_decap_8 FILLER_40_1142 ();
 sg13g2_decap_8 FILLER_40_1149 ();
 sg13g2_decap_8 FILLER_40_1156 ();
 sg13g2_decap_8 FILLER_40_1163 ();
 sg13g2_decap_8 FILLER_40_1170 ();
 sg13g2_decap_8 FILLER_40_1177 ();
 sg13g2_decap_8 FILLER_40_1184 ();
 sg13g2_decap_8 FILLER_40_1191 ();
 sg13g2_decap_8 FILLER_40_1198 ();
 sg13g2_decap_8 FILLER_40_1205 ();
 sg13g2_decap_8 FILLER_40_1212 ();
 sg13g2_decap_8 FILLER_40_1219 ();
 sg13g2_decap_8 FILLER_40_1226 ();
 sg13g2_decap_8 FILLER_40_1233 ();
 sg13g2_decap_8 FILLER_40_1240 ();
 sg13g2_decap_8 FILLER_40_1247 ();
 sg13g2_decap_8 FILLER_40_1254 ();
 sg13g2_decap_8 FILLER_40_1261 ();
 sg13g2_decap_8 FILLER_40_1268 ();
 sg13g2_decap_8 FILLER_40_1275 ();
 sg13g2_decap_8 FILLER_40_1282 ();
 sg13g2_decap_8 FILLER_40_1289 ();
 sg13g2_decap_8 FILLER_40_1296 ();
 sg13g2_decap_8 FILLER_40_1303 ();
 sg13g2_decap_4 FILLER_40_1310 ();
 sg13g2_fill_1 FILLER_40_1314 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_58 ();
 sg13g2_decap_4 FILLER_41_65 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_107 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_fill_1 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_decap_8 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_191 ();
 sg13g2_decap_8 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_4 FILLER_41_221 ();
 sg13g2_fill_2 FILLER_41_225 ();
 sg13g2_fill_2 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_423 ();
 sg13g2_fill_1 FILLER_41_427 ();
 sg13g2_fill_2 FILLER_41_436 ();
 sg13g2_decap_4 FILLER_41_452 ();
 sg13g2_fill_1 FILLER_41_456 ();
 sg13g2_decap_8 FILLER_41_461 ();
 sg13g2_fill_1 FILLER_41_468 ();
 sg13g2_decap_8 FILLER_41_487 ();
 sg13g2_decap_8 FILLER_41_494 ();
 sg13g2_fill_1 FILLER_41_501 ();
 sg13g2_fill_1 FILLER_41_510 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_decap_4 FILLER_41_535 ();
 sg13g2_fill_1 FILLER_41_544 ();
 sg13g2_fill_2 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_563 ();
 sg13g2_fill_1 FILLER_41_565 ();
 sg13g2_decap_4 FILLER_41_574 ();
 sg13g2_fill_2 FILLER_41_578 ();
 sg13g2_decap_4 FILLER_41_585 ();
 sg13g2_fill_1 FILLER_41_589 ();
 sg13g2_fill_2 FILLER_41_609 ();
 sg13g2_fill_1 FILLER_41_611 ();
 sg13g2_fill_1 FILLER_41_616 ();
 sg13g2_fill_2 FILLER_41_625 ();
 sg13g2_fill_2 FILLER_41_647 ();
 sg13g2_fill_1 FILLER_41_649 ();
 sg13g2_fill_1 FILLER_41_655 ();
 sg13g2_fill_2 FILLER_41_678 ();
 sg13g2_fill_1 FILLER_41_685 ();
 sg13g2_fill_2 FILLER_41_695 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_fill_1 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_fill_2 FILLER_41_728 ();
 sg13g2_fill_1 FILLER_41_787 ();
 sg13g2_decap_4 FILLER_41_793 ();
 sg13g2_fill_1 FILLER_41_797 ();
 sg13g2_fill_2 FILLER_41_802 ();
 sg13g2_fill_2 FILLER_41_840 ();
 sg13g2_fill_1 FILLER_41_842 ();
 sg13g2_decap_4 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_865 ();
 sg13g2_fill_1 FILLER_41_867 ();
 sg13g2_decap_4 FILLER_41_872 ();
 sg13g2_fill_2 FILLER_41_876 ();
 sg13g2_fill_2 FILLER_41_908 ();
 sg13g2_fill_1 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_954 ();
 sg13g2_fill_2 FILLER_41_969 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_fill_1 FILLER_41_996 ();
 sg13g2_fill_1 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1006 ();
 sg13g2_fill_1 FILLER_41_1013 ();
 sg13g2_fill_1 FILLER_41_1023 ();
 sg13g2_fill_2 FILLER_41_1029 ();
 sg13g2_fill_1 FILLER_41_1031 ();
 sg13g2_fill_2 FILLER_41_1045 ();
 sg13g2_decap_4 FILLER_41_1083 ();
 sg13g2_decap_8 FILLER_41_1097 ();
 sg13g2_fill_1 FILLER_41_1109 ();
 sg13g2_fill_1 FILLER_41_1114 ();
 sg13g2_decap_8 FILLER_41_1118 ();
 sg13g2_decap_8 FILLER_41_1125 ();
 sg13g2_decap_8 FILLER_41_1132 ();
 sg13g2_decap_8 FILLER_41_1139 ();
 sg13g2_decap_8 FILLER_41_1146 ();
 sg13g2_decap_8 FILLER_41_1153 ();
 sg13g2_decap_8 FILLER_41_1160 ();
 sg13g2_decap_8 FILLER_41_1167 ();
 sg13g2_decap_8 FILLER_41_1174 ();
 sg13g2_decap_8 FILLER_41_1181 ();
 sg13g2_decap_8 FILLER_41_1188 ();
 sg13g2_decap_8 FILLER_41_1195 ();
 sg13g2_decap_8 FILLER_41_1202 ();
 sg13g2_decap_8 FILLER_41_1209 ();
 sg13g2_decap_8 FILLER_41_1216 ();
 sg13g2_decap_8 FILLER_41_1223 ();
 sg13g2_decap_8 FILLER_41_1230 ();
 sg13g2_decap_8 FILLER_41_1237 ();
 sg13g2_decap_8 FILLER_41_1244 ();
 sg13g2_decap_8 FILLER_41_1251 ();
 sg13g2_decap_8 FILLER_41_1258 ();
 sg13g2_decap_8 FILLER_41_1265 ();
 sg13g2_decap_8 FILLER_41_1272 ();
 sg13g2_decap_8 FILLER_41_1279 ();
 sg13g2_decap_8 FILLER_41_1286 ();
 sg13g2_decap_8 FILLER_41_1293 ();
 sg13g2_decap_8 FILLER_41_1300 ();
 sg13g2_decap_8 FILLER_41_1307 ();
 sg13g2_fill_1 FILLER_41_1314 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_18 ();
 sg13g2_fill_2 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_44 ();
 sg13g2_fill_1 FILLER_42_53 ();
 sg13g2_decap_4 FILLER_42_80 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_fill_1 FILLER_42_181 ();
 sg13g2_fill_2 FILLER_42_229 ();
 sg13g2_fill_2 FILLER_42_262 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_269 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_1 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_283 ();
 sg13g2_decap_4 FILLER_42_290 ();
 sg13g2_fill_2 FILLER_42_294 ();
 sg13g2_fill_1 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_decap_4 FILLER_42_331 ();
 sg13g2_fill_2 FILLER_42_335 ();
 sg13g2_decap_8 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_362 ();
 sg13g2_decap_8 FILLER_42_369 ();
 sg13g2_decap_8 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_4 FILLER_42_400 ();
 sg13g2_fill_2 FILLER_42_404 ();
 sg13g2_decap_4 FILLER_42_421 ();
 sg13g2_fill_1 FILLER_42_430 ();
 sg13g2_fill_1 FILLER_42_438 ();
 sg13g2_decap_8 FILLER_42_447 ();
 sg13g2_fill_2 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_464 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_fill_2 FILLER_42_483 ();
 sg13g2_fill_1 FILLER_42_493 ();
 sg13g2_fill_2 FILLER_42_501 ();
 sg13g2_fill_1 FILLER_42_503 ();
 sg13g2_fill_2 FILLER_42_512 ();
 sg13g2_fill_1 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_551 ();
 sg13g2_fill_2 FILLER_42_574 ();
 sg13g2_fill_2 FILLER_42_594 ();
 sg13g2_fill_1 FILLER_42_612 ();
 sg13g2_decap_8 FILLER_42_622 ();
 sg13g2_fill_2 FILLER_42_629 ();
 sg13g2_fill_1 FILLER_42_631 ();
 sg13g2_fill_2 FILLER_42_645 ();
 sg13g2_fill_2 FILLER_42_673 ();
 sg13g2_decap_8 FILLER_42_688 ();
 sg13g2_fill_2 FILLER_42_704 ();
 sg13g2_fill_1 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_738 ();
 sg13g2_decap_8 FILLER_42_745 ();
 sg13g2_decap_4 FILLER_42_752 ();
 sg13g2_fill_1 FILLER_42_756 ();
 sg13g2_fill_1 FILLER_42_761 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_fill_2 FILLER_42_773 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_fill_1 FILLER_42_819 ();
 sg13g2_decap_4 FILLER_42_824 ();
 sg13g2_fill_2 FILLER_42_828 ();
 sg13g2_fill_1 FILLER_42_856 ();
 sg13g2_decap_4 FILLER_42_883 ();
 sg13g2_fill_2 FILLER_42_887 ();
 sg13g2_fill_1 FILLER_42_893 ();
 sg13g2_fill_1 FILLER_42_920 ();
 sg13g2_decap_8 FILLER_42_925 ();
 sg13g2_decap_8 FILLER_42_932 ();
 sg13g2_fill_2 FILLER_42_944 ();
 sg13g2_fill_2 FILLER_42_950 ();
 sg13g2_fill_1 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_1014 ();
 sg13g2_decap_4 FILLER_42_1043 ();
 sg13g2_fill_1 FILLER_42_1047 ();
 sg13g2_decap_4 FILLER_42_1053 ();
 sg13g2_fill_1 FILLER_42_1057 ();
 sg13g2_decap_8 FILLER_42_1062 ();
 sg13g2_fill_2 FILLER_42_1069 ();
 sg13g2_fill_2 FILLER_42_1097 ();
 sg13g2_fill_2 FILLER_42_1125 ();
 sg13g2_fill_1 FILLER_42_1127 ();
 sg13g2_decap_8 FILLER_42_1132 ();
 sg13g2_decap_8 FILLER_42_1139 ();
 sg13g2_decap_8 FILLER_42_1146 ();
 sg13g2_decap_8 FILLER_42_1153 ();
 sg13g2_decap_8 FILLER_42_1160 ();
 sg13g2_decap_8 FILLER_42_1167 ();
 sg13g2_decap_8 FILLER_42_1174 ();
 sg13g2_decap_8 FILLER_42_1181 ();
 sg13g2_decap_8 FILLER_42_1188 ();
 sg13g2_decap_8 FILLER_42_1195 ();
 sg13g2_decap_8 FILLER_42_1202 ();
 sg13g2_decap_8 FILLER_42_1209 ();
 sg13g2_decap_8 FILLER_42_1216 ();
 sg13g2_decap_8 FILLER_42_1223 ();
 sg13g2_decap_8 FILLER_42_1230 ();
 sg13g2_decap_8 FILLER_42_1237 ();
 sg13g2_decap_8 FILLER_42_1244 ();
 sg13g2_decap_8 FILLER_42_1251 ();
 sg13g2_decap_8 FILLER_42_1258 ();
 sg13g2_decap_8 FILLER_42_1265 ();
 sg13g2_decap_8 FILLER_42_1272 ();
 sg13g2_decap_8 FILLER_42_1279 ();
 sg13g2_decap_8 FILLER_42_1286 ();
 sg13g2_decap_8 FILLER_42_1293 ();
 sg13g2_decap_8 FILLER_42_1300 ();
 sg13g2_decap_8 FILLER_42_1307 ();
 sg13g2_fill_1 FILLER_42_1314 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_41 ();
 sg13g2_fill_2 FILLER_43_48 ();
 sg13g2_decap_4 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_2 FILLER_43_64 ();
 sg13g2_fill_1 FILLER_43_66 ();
 sg13g2_decap_8 FILLER_43_72 ();
 sg13g2_decap_8 FILLER_43_79 ();
 sg13g2_decap_8 FILLER_43_86 ();
 sg13g2_decap_4 FILLER_43_93 ();
 sg13g2_decap_8 FILLER_43_101 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_decap_4 FILLER_43_115 ();
 sg13g2_fill_2 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_125 ();
 sg13g2_decap_8 FILLER_43_132 ();
 sg13g2_decap_8 FILLER_43_139 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_158 ();
 sg13g2_fill_2 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_decap_4 FILLER_43_187 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_fill_2 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_205 ();
 sg13g2_fill_2 FILLER_43_214 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_246 ();
 sg13g2_fill_2 FILLER_43_253 ();
 sg13g2_fill_1 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_266 ();
 sg13g2_fill_2 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_363 ();
 sg13g2_decap_4 FILLER_43_370 ();
 sg13g2_fill_2 FILLER_43_401 ();
 sg13g2_decap_4 FILLER_43_410 ();
 sg13g2_fill_2 FILLER_43_448 ();
 sg13g2_fill_1 FILLER_43_450 ();
 sg13g2_fill_2 FILLER_43_461 ();
 sg13g2_decap_8 FILLER_43_482 ();
 sg13g2_decap_4 FILLER_43_489 ();
 sg13g2_fill_2 FILLER_43_493 ();
 sg13g2_fill_2 FILLER_43_536 ();
 sg13g2_fill_1 FILLER_43_538 ();
 sg13g2_fill_2 FILLER_43_562 ();
 sg13g2_fill_2 FILLER_43_569 ();
 sg13g2_decap_8 FILLER_43_585 ();
 sg13g2_fill_2 FILLER_43_592 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_fill_1 FILLER_43_600 ();
 sg13g2_fill_2 FILLER_43_606 ();
 sg13g2_fill_1 FILLER_43_608 ();
 sg13g2_fill_2 FILLER_43_619 ();
 sg13g2_fill_2 FILLER_43_642 ();
 sg13g2_fill_1 FILLER_43_644 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_decap_4 FILLER_43_671 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_fill_2 FILLER_43_686 ();
 sg13g2_fill_2 FILLER_43_694 ();
 sg13g2_fill_2 FILLER_43_711 ();
 sg13g2_fill_1 FILLER_43_724 ();
 sg13g2_fill_2 FILLER_43_754 ();
 sg13g2_decap_4 FILLER_43_782 ();
 sg13g2_fill_2 FILLER_43_811 ();
 sg13g2_fill_1 FILLER_43_813 ();
 sg13g2_fill_2 FILLER_43_822 ();
 sg13g2_fill_1 FILLER_43_824 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_fill_1 FILLER_43_836 ();
 sg13g2_decap_4 FILLER_43_862 ();
 sg13g2_fill_2 FILLER_43_866 ();
 sg13g2_fill_2 FILLER_43_872 ();
 sg13g2_fill_1 FILLER_43_878 ();
 sg13g2_fill_2 FILLER_43_888 ();
 sg13g2_fill_1 FILLER_43_895 ();
 sg13g2_decap_4 FILLER_43_901 ();
 sg13g2_fill_2 FILLER_43_913 ();
 sg13g2_fill_1 FILLER_43_915 ();
 sg13g2_fill_2 FILLER_43_921 ();
 sg13g2_decap_4 FILLER_43_932 ();
 sg13g2_fill_1 FILLER_43_962 ();
 sg13g2_decap_4 FILLER_43_1003 ();
 sg13g2_fill_1 FILLER_43_1007 ();
 sg13g2_fill_2 FILLER_43_1075 ();
 sg13g2_fill_1 FILLER_43_1086 ();
 sg13g2_decap_4 FILLER_43_1090 ();
 sg13g2_fill_2 FILLER_43_1104 ();
 sg13g2_fill_1 FILLER_43_1106 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1178 ();
 sg13g2_decap_8 FILLER_43_1185 ();
 sg13g2_decap_8 FILLER_43_1192 ();
 sg13g2_decap_8 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_decap_8 FILLER_43_1213 ();
 sg13g2_decap_8 FILLER_43_1220 ();
 sg13g2_decap_8 FILLER_43_1227 ();
 sg13g2_decap_8 FILLER_43_1234 ();
 sg13g2_decap_8 FILLER_43_1241 ();
 sg13g2_decap_8 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1255 ();
 sg13g2_decap_8 FILLER_43_1262 ();
 sg13g2_decap_8 FILLER_43_1269 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_4 FILLER_43_1311 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_27 ();
 sg13g2_decap_4 FILLER_44_34 ();
 sg13g2_fill_2 FILLER_44_54 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_decap_4 FILLER_44_83 ();
 sg13g2_fill_1 FILLER_44_87 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_103 ();
 sg13g2_fill_1 FILLER_44_105 ();
 sg13g2_fill_2 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_fill_1 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_219 ();
 sg13g2_fill_2 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_fill_2 FILLER_44_337 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_2 FILLER_44_385 ();
 sg13g2_decap_4 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_448 ();
 sg13g2_fill_1 FILLER_44_450 ();
 sg13g2_fill_1 FILLER_44_485 ();
 sg13g2_fill_1 FILLER_44_509 ();
 sg13g2_decap_4 FILLER_44_515 ();
 sg13g2_fill_2 FILLER_44_519 ();
 sg13g2_decap_4 FILLER_44_531 ();
 sg13g2_decap_8 FILLER_44_544 ();
 sg13g2_decap_8 FILLER_44_551 ();
 sg13g2_fill_2 FILLER_44_572 ();
 sg13g2_decap_4 FILLER_44_580 ();
 sg13g2_fill_2 FILLER_44_605 ();
 sg13g2_decap_8 FILLER_44_619 ();
 sg13g2_fill_1 FILLER_44_626 ();
 sg13g2_decap_4 FILLER_44_646 ();
 sg13g2_fill_1 FILLER_44_650 ();
 sg13g2_fill_2 FILLER_44_661 ();
 sg13g2_fill_2 FILLER_44_672 ();
 sg13g2_fill_2 FILLER_44_688 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_fill_2 FILLER_44_700 ();
 sg13g2_decap_4 FILLER_44_706 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_fill_1 FILLER_44_740 ();
 sg13g2_decap_8 FILLER_44_759 ();
 sg13g2_fill_1 FILLER_44_766 ();
 sg13g2_decap_4 FILLER_44_771 ();
 sg13g2_fill_2 FILLER_44_775 ();
 sg13g2_fill_2 FILLER_44_786 ();
 sg13g2_fill_2 FILLER_44_809 ();
 sg13g2_fill_2 FILLER_44_837 ();
 sg13g2_fill_1 FILLER_44_839 ();
 sg13g2_fill_2 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_44_873 ();
 sg13g2_fill_1 FILLER_44_875 ();
 sg13g2_decap_4 FILLER_44_907 ();
 sg13g2_fill_1 FILLER_44_911 ();
 sg13g2_decap_4 FILLER_44_945 ();
 sg13g2_fill_1 FILLER_44_949 ();
 sg13g2_decap_8 FILLER_44_961 ();
 sg13g2_decap_8 FILLER_44_968 ();
 sg13g2_decap_8 FILLER_44_975 ();
 sg13g2_fill_2 FILLER_44_982 ();
 sg13g2_fill_1 FILLER_44_988 ();
 sg13g2_fill_1 FILLER_44_1018 ();
 sg13g2_decap_8 FILLER_44_1023 ();
 sg13g2_fill_1 FILLER_44_1034 ();
 sg13g2_decap_8 FILLER_44_1040 ();
 sg13g2_fill_1 FILLER_44_1047 ();
 sg13g2_fill_1 FILLER_44_1060 ();
 sg13g2_fill_2 FILLER_44_1065 ();
 sg13g2_fill_1 FILLER_44_1067 ();
 sg13g2_decap_8 FILLER_44_1104 ();
 sg13g2_fill_1 FILLER_44_1111 ();
 sg13g2_decap_8 FILLER_44_1138 ();
 sg13g2_decap_8 FILLER_44_1145 ();
 sg13g2_decap_8 FILLER_44_1152 ();
 sg13g2_decap_8 FILLER_44_1159 ();
 sg13g2_decap_8 FILLER_44_1166 ();
 sg13g2_decap_8 FILLER_44_1173 ();
 sg13g2_decap_8 FILLER_44_1180 ();
 sg13g2_decap_8 FILLER_44_1187 ();
 sg13g2_decap_8 FILLER_44_1194 ();
 sg13g2_decap_8 FILLER_44_1201 ();
 sg13g2_decap_8 FILLER_44_1208 ();
 sg13g2_decap_8 FILLER_44_1215 ();
 sg13g2_decap_8 FILLER_44_1222 ();
 sg13g2_decap_8 FILLER_44_1229 ();
 sg13g2_decap_8 FILLER_44_1236 ();
 sg13g2_decap_8 FILLER_44_1243 ();
 sg13g2_decap_8 FILLER_44_1250 ();
 sg13g2_decap_8 FILLER_44_1257 ();
 sg13g2_decap_8 FILLER_44_1264 ();
 sg13g2_decap_8 FILLER_44_1271 ();
 sg13g2_decap_8 FILLER_44_1278 ();
 sg13g2_decap_8 FILLER_44_1285 ();
 sg13g2_decap_8 FILLER_44_1292 ();
 sg13g2_decap_8 FILLER_44_1299 ();
 sg13g2_decap_8 FILLER_44_1306 ();
 sg13g2_fill_2 FILLER_44_1313 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_decap_4 FILLER_45_16 ();
 sg13g2_fill_1 FILLER_45_24 ();
 sg13g2_fill_2 FILLER_45_70 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_decap_8 FILLER_45_135 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_decap_8 FILLER_45_169 ();
 sg13g2_decap_8 FILLER_45_176 ();
 sg13g2_fill_2 FILLER_45_183 ();
 sg13g2_fill_1 FILLER_45_185 ();
 sg13g2_decap_4 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_4 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_239 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_fill_1 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_fill_1 FILLER_45_314 ();
 sg13g2_decap_4 FILLER_45_323 ();
 sg13g2_fill_1 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_fill_2 FILLER_45_356 ();
 sg13g2_decap_8 FILLER_45_362 ();
 sg13g2_decap_4 FILLER_45_369 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_decap_4 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_407 ();
 sg13g2_fill_1 FILLER_45_414 ();
 sg13g2_decap_8 FILLER_45_421 ();
 sg13g2_decap_8 FILLER_45_428 ();
 sg13g2_fill_2 FILLER_45_435 ();
 sg13g2_fill_1 FILLER_45_437 ();
 sg13g2_fill_2 FILLER_45_464 ();
 sg13g2_fill_1 FILLER_45_466 ();
 sg13g2_decap_4 FILLER_45_476 ();
 sg13g2_fill_2 FILLER_45_506 ();
 sg13g2_decap_4 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_2 FILLER_45_540 ();
 sg13g2_decap_4 FILLER_45_550 ();
 sg13g2_fill_1 FILLER_45_563 ();
 sg13g2_fill_2 FILLER_45_572 ();
 sg13g2_fill_1 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_586 ();
 sg13g2_decap_4 FILLER_45_593 ();
 sg13g2_fill_1 FILLER_45_597 ();
 sg13g2_decap_8 FILLER_45_613 ();
 sg13g2_fill_2 FILLER_45_620 ();
 sg13g2_decap_4 FILLER_45_636 ();
 sg13g2_decap_4 FILLER_45_663 ();
 sg13g2_fill_1 FILLER_45_672 ();
 sg13g2_fill_2 FILLER_45_691 ();
 sg13g2_fill_1 FILLER_45_693 ();
 sg13g2_fill_1 FILLER_45_704 ();
 sg13g2_fill_1 FILLER_45_713 ();
 sg13g2_decap_4 FILLER_45_719 ();
 sg13g2_decap_4 FILLER_45_727 ();
 sg13g2_decap_8 FILLER_45_744 ();
 sg13g2_decap_4 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_4 FILLER_45_766 ();
 sg13g2_fill_2 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_832 ();
 sg13g2_decap_8 FILLER_45_839 ();
 sg13g2_decap_8 FILLER_45_846 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_fill_1 FILLER_45_860 ();
 sg13g2_fill_2 FILLER_45_869 ();
 sg13g2_fill_2 FILLER_45_875 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_decap_8 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_895 ();
 sg13g2_decap_4 FILLER_45_919 ();
 sg13g2_fill_2 FILLER_45_923 ();
 sg13g2_fill_1 FILLER_45_935 ();
 sg13g2_fill_2 FILLER_45_962 ();
 sg13g2_fill_1 FILLER_45_964 ();
 sg13g2_fill_2 FILLER_45_1025 ();
 sg13g2_fill_1 FILLER_45_1027 ();
 sg13g2_decap_8 FILLER_45_1074 ();
 sg13g2_decap_4 FILLER_45_1099 ();
 sg13g2_fill_2 FILLER_45_1130 ();
 sg13g2_fill_1 FILLER_45_1132 ();
 sg13g2_decap_8 FILLER_45_1136 ();
 sg13g2_decap_8 FILLER_45_1143 ();
 sg13g2_decap_8 FILLER_45_1150 ();
 sg13g2_decap_8 FILLER_45_1157 ();
 sg13g2_decap_8 FILLER_45_1164 ();
 sg13g2_decap_8 FILLER_45_1171 ();
 sg13g2_decap_8 FILLER_45_1178 ();
 sg13g2_decap_8 FILLER_45_1185 ();
 sg13g2_decap_8 FILLER_45_1192 ();
 sg13g2_decap_8 FILLER_45_1199 ();
 sg13g2_decap_8 FILLER_45_1206 ();
 sg13g2_decap_8 FILLER_45_1213 ();
 sg13g2_decap_8 FILLER_45_1220 ();
 sg13g2_decap_8 FILLER_45_1227 ();
 sg13g2_decap_8 FILLER_45_1234 ();
 sg13g2_decap_8 FILLER_45_1241 ();
 sg13g2_decap_8 FILLER_45_1248 ();
 sg13g2_decap_8 FILLER_45_1255 ();
 sg13g2_decap_8 FILLER_45_1262 ();
 sg13g2_decap_8 FILLER_45_1269 ();
 sg13g2_decap_8 FILLER_45_1276 ();
 sg13g2_decap_8 FILLER_45_1283 ();
 sg13g2_decap_8 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1297 ();
 sg13g2_decap_8 FILLER_45_1304 ();
 sg13g2_decap_4 FILLER_45_1311 ();
 sg13g2_decap_8 FILLER_46_39 ();
 sg13g2_fill_1 FILLER_46_55 ();
 sg13g2_decap_8 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_68 ();
 sg13g2_decap_4 FILLER_46_75 ();
 sg13g2_fill_2 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_94 ();
 sg13g2_fill_2 FILLER_46_124 ();
 sg13g2_decap_4 FILLER_46_191 ();
 sg13g2_fill_2 FILLER_46_206 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_decap_8 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_decap_4 FILLER_46_241 ();
 sg13g2_fill_1 FILLER_46_245 ();
 sg13g2_fill_2 FILLER_46_272 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_281 ();
 sg13g2_fill_2 FILLER_46_296 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_345 ();
 sg13g2_fill_1 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_420 ();
 sg13g2_fill_1 FILLER_46_422 ();
 sg13g2_decap_4 FILLER_46_428 ();
 sg13g2_fill_1 FILLER_46_432 ();
 sg13g2_fill_2 FILLER_46_437 ();
 sg13g2_decap_8 FILLER_46_456 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_decap_4 FILLER_46_482 ();
 sg13g2_fill_2 FILLER_46_486 ();
 sg13g2_fill_1 FILLER_46_494 ();
 sg13g2_fill_2 FILLER_46_504 ();
 sg13g2_fill_1 FILLER_46_506 ();
 sg13g2_fill_1 FILLER_46_511 ();
 sg13g2_fill_2 FILLER_46_540 ();
 sg13g2_fill_2 FILLER_46_553 ();
 sg13g2_fill_1 FILLER_46_560 ();
 sg13g2_fill_2 FILLER_46_570 ();
 sg13g2_fill_1 FILLER_46_591 ();
 sg13g2_fill_2 FILLER_46_611 ();
 sg13g2_fill_1 FILLER_46_613 ();
 sg13g2_decap_4 FILLER_46_618 ();
 sg13g2_fill_1 FILLER_46_641 ();
 sg13g2_fill_2 FILLER_46_657 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_fill_2 FILLER_46_675 ();
 sg13g2_fill_1 FILLER_46_677 ();
 sg13g2_fill_2 FILLER_46_689 ();
 sg13g2_decap_4 FILLER_46_705 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_decap_4 FILLER_46_715 ();
 sg13g2_fill_2 FILLER_46_731 ();
 sg13g2_fill_1 FILLER_46_733 ();
 sg13g2_decap_8 FILLER_46_810 ();
 sg13g2_fill_2 FILLER_46_817 ();
 sg13g2_fill_1 FILLER_46_819 ();
 sg13g2_decap_4 FILLER_46_855 ();
 sg13g2_fill_2 FILLER_46_864 ();
 sg13g2_fill_1 FILLER_46_866 ();
 sg13g2_fill_1 FILLER_46_875 ();
 sg13g2_fill_1 FILLER_46_910 ();
 sg13g2_decap_4 FILLER_46_916 ();
 sg13g2_fill_2 FILLER_46_920 ();
 sg13g2_decap_8 FILLER_46_934 ();
 sg13g2_fill_2 FILLER_46_941 ();
 sg13g2_fill_2 FILLER_46_960 ();
 sg13g2_decap_8 FILLER_46_984 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_998 ();
 sg13g2_decap_4 FILLER_46_1005 ();
 sg13g2_fill_1 FILLER_46_1009 ();
 sg13g2_fill_2 FILLER_46_1018 ();
 sg13g2_fill_1 FILLER_46_1020 ();
 sg13g2_decap_4 FILLER_46_1026 ();
 sg13g2_fill_2 FILLER_46_1030 ();
 sg13g2_decap_8 FILLER_46_1041 ();
 sg13g2_fill_1 FILLER_46_1048 ();
 sg13g2_fill_2 FILLER_46_1059 ();
 sg13g2_fill_1 FILLER_46_1061 ();
 sg13g2_fill_2 FILLER_46_1081 ();
 sg13g2_decap_4 FILLER_46_1113 ();
 sg13g2_fill_1 FILLER_46_1117 ();
 sg13g2_decap_8 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_decap_8 FILLER_46_1158 ();
 sg13g2_decap_8 FILLER_46_1165 ();
 sg13g2_decap_8 FILLER_46_1172 ();
 sg13g2_decap_8 FILLER_46_1179 ();
 sg13g2_decap_8 FILLER_46_1186 ();
 sg13g2_decap_8 FILLER_46_1193 ();
 sg13g2_decap_8 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1207 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_decap_8 FILLER_46_1221 ();
 sg13g2_decap_8 FILLER_46_1228 ();
 sg13g2_decap_8 FILLER_46_1235 ();
 sg13g2_decap_8 FILLER_46_1242 ();
 sg13g2_decap_8 FILLER_46_1249 ();
 sg13g2_decap_8 FILLER_46_1256 ();
 sg13g2_decap_8 FILLER_46_1263 ();
 sg13g2_decap_8 FILLER_46_1270 ();
 sg13g2_decap_8 FILLER_46_1277 ();
 sg13g2_decap_8 FILLER_46_1284 ();
 sg13g2_decap_8 FILLER_46_1291 ();
 sg13g2_decap_8 FILLER_46_1298 ();
 sg13g2_decap_8 FILLER_46_1305 ();
 sg13g2_fill_2 FILLER_46_1312 ();
 sg13g2_fill_1 FILLER_46_1314 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_decap_8 FILLER_47_143 ();
 sg13g2_decap_4 FILLER_47_150 ();
 sg13g2_fill_2 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_fill_1 FILLER_47_203 ();
 sg13g2_decap_4 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_fill_2 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_fill_2 FILLER_47_422 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_4 FILLER_47_446 ();
 sg13g2_fill_2 FILLER_47_450 ();
 sg13g2_decap_8 FILLER_47_465 ();
 sg13g2_decap_4 FILLER_47_472 ();
 sg13g2_fill_2 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_484 ();
 sg13g2_decap_8 FILLER_47_491 ();
 sg13g2_fill_1 FILLER_47_498 ();
 sg13g2_decap_4 FILLER_47_522 ();
 sg13g2_fill_2 FILLER_47_526 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_fill_2 FILLER_47_551 ();
 sg13g2_fill_2 FILLER_47_568 ();
 sg13g2_fill_2 FILLER_47_579 ();
 sg13g2_fill_1 FILLER_47_589 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_fill_1 FILLER_47_602 ();
 sg13g2_fill_1 FILLER_47_627 ();
 sg13g2_decap_8 FILLER_47_641 ();
 sg13g2_fill_1 FILLER_47_648 ();
 sg13g2_fill_1 FILLER_47_653 ();
 sg13g2_fill_2 FILLER_47_671 ();
 sg13g2_fill_2 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_679 ();
 sg13g2_fill_2 FILLER_47_693 ();
 sg13g2_fill_1 FILLER_47_695 ();
 sg13g2_fill_2 FILLER_47_718 ();
 sg13g2_decap_4 FILLER_47_736 ();
 sg13g2_fill_2 FILLER_47_740 ();
 sg13g2_decap_4 FILLER_47_769 ();
 sg13g2_fill_2 FILLER_47_773 ();
 sg13g2_decap_4 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_793 ();
 sg13g2_decap_8 FILLER_47_816 ();
 sg13g2_fill_1 FILLER_47_823 ();
 sg13g2_fill_2 FILLER_47_858 ();
 sg13g2_fill_1 FILLER_47_860 ();
 sg13g2_fill_2 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_47_891 ();
 sg13g2_fill_1 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_912 ();
 sg13g2_fill_1 FILLER_47_919 ();
 sg13g2_fill_2 FILLER_47_925 ();
 sg13g2_fill_2 FILLER_47_943 ();
 sg13g2_fill_1 FILLER_47_945 ();
 sg13g2_fill_2 FILLER_47_954 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_fill_2 FILLER_47_1017 ();
 sg13g2_fill_1 FILLER_47_1032 ();
 sg13g2_decap_4 FILLER_47_1041 ();
 sg13g2_decap_4 FILLER_47_1068 ();
 sg13g2_fill_1 FILLER_47_1077 ();
 sg13g2_decap_8 FILLER_47_1119 ();
 sg13g2_fill_2 FILLER_47_1126 ();
 sg13g2_fill_1 FILLER_47_1128 ();
 sg13g2_decap_8 FILLER_47_1133 ();
 sg13g2_decap_8 FILLER_47_1140 ();
 sg13g2_decap_8 FILLER_47_1147 ();
 sg13g2_decap_8 FILLER_47_1154 ();
 sg13g2_decap_8 FILLER_47_1161 ();
 sg13g2_decap_8 FILLER_47_1168 ();
 sg13g2_decap_8 FILLER_47_1175 ();
 sg13g2_decap_8 FILLER_47_1182 ();
 sg13g2_decap_8 FILLER_47_1189 ();
 sg13g2_decap_8 FILLER_47_1196 ();
 sg13g2_decap_8 FILLER_47_1203 ();
 sg13g2_decap_8 FILLER_47_1210 ();
 sg13g2_decap_8 FILLER_47_1217 ();
 sg13g2_decap_8 FILLER_47_1224 ();
 sg13g2_decap_8 FILLER_47_1231 ();
 sg13g2_decap_8 FILLER_47_1238 ();
 sg13g2_decap_8 FILLER_47_1245 ();
 sg13g2_decap_8 FILLER_47_1252 ();
 sg13g2_decap_8 FILLER_47_1259 ();
 sg13g2_decap_8 FILLER_47_1266 ();
 sg13g2_decap_8 FILLER_47_1273 ();
 sg13g2_decap_8 FILLER_47_1280 ();
 sg13g2_decap_8 FILLER_47_1287 ();
 sg13g2_decap_8 FILLER_47_1294 ();
 sg13g2_decap_8 FILLER_47_1301 ();
 sg13g2_decap_8 FILLER_47_1308 ();
 sg13g2_decap_4 FILLER_48_62 ();
 sg13g2_decap_4 FILLER_48_92 ();
 sg13g2_fill_2 FILLER_48_96 ();
 sg13g2_fill_2 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_108 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_decap_4 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_132 ();
 sg13g2_fill_1 FILLER_48_134 ();
 sg13g2_decap_8 FILLER_48_162 ();
 sg13g2_decap_8 FILLER_48_169 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_decap_8 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_190 ();
 sg13g2_fill_1 FILLER_48_192 ();
 sg13g2_decap_4 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_246 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_2 FILLER_48_284 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_1 FILLER_48_297 ();
 sg13g2_decap_4 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_decap_4 FILLER_48_386 ();
 sg13g2_fill_1 FILLER_48_390 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_decap_8 FILLER_48_454 ();
 sg13g2_fill_2 FILLER_48_471 ();
 sg13g2_decap_4 FILLER_48_524 ();
 sg13g2_decap_4 FILLER_48_542 ();
 sg13g2_fill_1 FILLER_48_546 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_fill_2 FILLER_48_581 ();
 sg13g2_fill_1 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_605 ();
 sg13g2_fill_2 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_fill_1 FILLER_48_652 ();
 sg13g2_fill_1 FILLER_48_665 ();
 sg13g2_fill_2 FILLER_48_671 ();
 sg13g2_fill_1 FILLER_48_673 ();
 sg13g2_decap_4 FILLER_48_687 ();
 sg13g2_fill_2 FILLER_48_691 ();
 sg13g2_decap_8 FILLER_48_706 ();
 sg13g2_decap_8 FILLER_48_713 ();
 sg13g2_fill_1 FILLER_48_732 ();
 sg13g2_decap_4 FILLER_48_746 ();
 sg13g2_fill_1 FILLER_48_750 ();
 sg13g2_decap_4 FILLER_48_790 ();
 sg13g2_decap_4 FILLER_48_833 ();
 sg13g2_fill_1 FILLER_48_837 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_fill_2 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_fill_1 FILLER_48_877 ();
 sg13g2_fill_2 FILLER_48_904 ();
 sg13g2_decap_8 FILLER_48_932 ();
 sg13g2_fill_2 FILLER_48_939 ();
 sg13g2_decap_8 FILLER_48_946 ();
 sg13g2_decap_8 FILLER_48_969 ();
 sg13g2_fill_1 FILLER_48_976 ();
 sg13g2_decap_8 FILLER_48_986 ();
 sg13g2_decap_4 FILLER_48_993 ();
 sg13g2_decap_8 FILLER_48_1013 ();
 sg13g2_decap_8 FILLER_48_1020 ();
 sg13g2_fill_2 FILLER_48_1027 ();
 sg13g2_fill_1 FILLER_48_1029 ();
 sg13g2_fill_2 FILLER_48_1035 ();
 sg13g2_decap_8 FILLER_48_1042 ();
 sg13g2_fill_2 FILLER_48_1049 ();
 sg13g2_decap_4 FILLER_48_1075 ();
 sg13g2_fill_1 FILLER_48_1079 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_4 FILLER_48_1099 ();
 sg13g2_fill_1 FILLER_48_1103 ();
 sg13g2_decap_4 FILLER_48_1109 ();
 sg13g2_decap_8 FILLER_48_1121 ();
 sg13g2_decap_8 FILLER_48_1128 ();
 sg13g2_decap_8 FILLER_48_1135 ();
 sg13g2_decap_8 FILLER_48_1142 ();
 sg13g2_decap_8 FILLER_48_1149 ();
 sg13g2_decap_8 FILLER_48_1156 ();
 sg13g2_decap_8 FILLER_48_1163 ();
 sg13g2_decap_8 FILLER_48_1170 ();
 sg13g2_decap_8 FILLER_48_1177 ();
 sg13g2_decap_8 FILLER_48_1184 ();
 sg13g2_decap_8 FILLER_48_1191 ();
 sg13g2_decap_8 FILLER_48_1198 ();
 sg13g2_decap_8 FILLER_48_1205 ();
 sg13g2_decap_8 FILLER_48_1212 ();
 sg13g2_decap_8 FILLER_48_1219 ();
 sg13g2_decap_8 FILLER_48_1226 ();
 sg13g2_decap_8 FILLER_48_1233 ();
 sg13g2_decap_8 FILLER_48_1240 ();
 sg13g2_decap_8 FILLER_48_1247 ();
 sg13g2_decap_8 FILLER_48_1254 ();
 sg13g2_decap_8 FILLER_48_1261 ();
 sg13g2_decap_8 FILLER_48_1268 ();
 sg13g2_decap_8 FILLER_48_1275 ();
 sg13g2_decap_8 FILLER_48_1282 ();
 sg13g2_decap_8 FILLER_48_1289 ();
 sg13g2_decap_8 FILLER_48_1296 ();
 sg13g2_decap_8 FILLER_48_1303 ();
 sg13g2_decap_4 FILLER_48_1310 ();
 sg13g2_fill_1 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_49_30 ();
 sg13g2_decap_4 FILLER_49_37 ();
 sg13g2_fill_2 FILLER_49_41 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_decap_8 FILLER_49_69 ();
 sg13g2_fill_2 FILLER_49_76 ();
 sg13g2_decap_4 FILLER_49_86 ();
 sg13g2_decap_4 FILLER_49_94 ();
 sg13g2_decap_4 FILLER_49_136 ();
 sg13g2_fill_1 FILLER_49_140 ();
 sg13g2_fill_2 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_197 ();
 sg13g2_fill_2 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_216 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_decap_4 FILLER_49_237 ();
 sg13g2_decap_4 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_decap_4 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_338 ();
 sg13g2_fill_2 FILLER_49_342 ();
 sg13g2_fill_2 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_fill_2 FILLER_49_366 ();
 sg13g2_fill_2 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_414 ();
 sg13g2_fill_1 FILLER_49_416 ();
 sg13g2_fill_2 FILLER_49_427 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_decap_4 FILLER_49_435 ();
 sg13g2_fill_1 FILLER_49_439 ();
 sg13g2_fill_2 FILLER_49_450 ();
 sg13g2_fill_2 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_492 ();
 sg13g2_decap_4 FILLER_49_499 ();
 sg13g2_fill_2 FILLER_49_515 ();
 sg13g2_fill_2 FILLER_49_523 ();
 sg13g2_decap_4 FILLER_49_529 ();
 sg13g2_fill_2 FILLER_49_533 ();
 sg13g2_fill_1 FILLER_49_550 ();
 sg13g2_decap_4 FILLER_49_571 ();
 sg13g2_fill_2 FILLER_49_575 ();
 sg13g2_fill_2 FILLER_49_582 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_fill_1 FILLER_49_595 ();
 sg13g2_fill_1 FILLER_49_619 ();
 sg13g2_decap_8 FILLER_49_634 ();
 sg13g2_decap_4 FILLER_49_641 ();
 sg13g2_fill_2 FILLER_49_645 ();
 sg13g2_decap_4 FILLER_49_651 ();
 sg13g2_fill_2 FILLER_49_671 ();
 sg13g2_fill_1 FILLER_49_673 ();
 sg13g2_decap_8 FILLER_49_688 ();
 sg13g2_fill_2 FILLER_49_728 ();
 sg13g2_fill_1 FILLER_49_730 ();
 sg13g2_decap_8 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_804 ();
 sg13g2_fill_2 FILLER_49_811 ();
 sg13g2_fill_2 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_fill_1 FILLER_49_846 ();
 sg13g2_fill_2 FILLER_49_867 ();
 sg13g2_fill_2 FILLER_49_874 ();
 sg13g2_fill_2 FILLER_49_880 ();
 sg13g2_fill_1 FILLER_49_887 ();
 sg13g2_decap_8 FILLER_49_892 ();
 sg13g2_decap_8 FILLER_49_899 ();
 sg13g2_fill_1 FILLER_49_906 ();
 sg13g2_fill_1 FILLER_49_912 ();
 sg13g2_fill_1 FILLER_49_925 ();
 sg13g2_fill_1 FILLER_49_956 ();
 sg13g2_decap_4 FILLER_49_966 ();
 sg13g2_fill_2 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_998 ();
 sg13g2_fill_1 FILLER_49_1000 ();
 sg13g2_fill_2 FILLER_49_1032 ();
 sg13g2_fill_1 FILLER_49_1034 ();
 sg13g2_fill_1 FILLER_49_1050 ();
 sg13g2_fill_1 FILLER_49_1056 ();
 sg13g2_decap_4 FILLER_49_1070 ();
 sg13g2_fill_2 FILLER_49_1074 ();
 sg13g2_fill_1 FILLER_49_1102 ();
 sg13g2_decap_8 FILLER_49_1132 ();
 sg13g2_decap_8 FILLER_49_1139 ();
 sg13g2_decap_8 FILLER_49_1146 ();
 sg13g2_decap_8 FILLER_49_1153 ();
 sg13g2_decap_8 FILLER_49_1160 ();
 sg13g2_decap_8 FILLER_49_1167 ();
 sg13g2_decap_8 FILLER_49_1174 ();
 sg13g2_decap_8 FILLER_49_1181 ();
 sg13g2_decap_8 FILLER_49_1188 ();
 sg13g2_decap_8 FILLER_49_1195 ();
 sg13g2_decap_8 FILLER_49_1202 ();
 sg13g2_decap_8 FILLER_49_1209 ();
 sg13g2_decap_8 FILLER_49_1216 ();
 sg13g2_decap_8 FILLER_49_1223 ();
 sg13g2_decap_8 FILLER_49_1230 ();
 sg13g2_decap_8 FILLER_49_1237 ();
 sg13g2_decap_8 FILLER_49_1244 ();
 sg13g2_decap_8 FILLER_49_1251 ();
 sg13g2_decap_8 FILLER_49_1258 ();
 sg13g2_decap_8 FILLER_49_1265 ();
 sg13g2_decap_8 FILLER_49_1272 ();
 sg13g2_decap_8 FILLER_49_1279 ();
 sg13g2_decap_8 FILLER_49_1286 ();
 sg13g2_decap_8 FILLER_49_1293 ();
 sg13g2_decap_8 FILLER_49_1300 ();
 sg13g2_decap_8 FILLER_49_1307 ();
 sg13g2_fill_1 FILLER_49_1314 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_30 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_decap_4 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_decap_4 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_decap_8 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_188 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_233 ();
 sg13g2_fill_2 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_259 ();
 sg13g2_fill_1 FILLER_50_261 ();
 sg13g2_fill_2 FILLER_50_297 ();
 sg13g2_fill_1 FILLER_50_299 ();
 sg13g2_decap_8 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_349 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_fill_1 FILLER_50_394 ();
 sg13g2_fill_2 FILLER_50_410 ();
 sg13g2_fill_1 FILLER_50_412 ();
 sg13g2_decap_4 FILLER_50_418 ();
 sg13g2_decap_4 FILLER_50_430 ();
 sg13g2_decap_8 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_fill_2 FILLER_50_459 ();
 sg13g2_fill_1 FILLER_50_466 ();
 sg13g2_decap_4 FILLER_50_482 ();
 sg13g2_fill_2 FILLER_50_500 ();
 sg13g2_fill_1 FILLER_50_502 ();
 sg13g2_fill_2 FILLER_50_521 ();
 sg13g2_decap_8 FILLER_50_543 ();
 sg13g2_fill_2 FILLER_50_550 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_decap_8 FILLER_50_606 ();
 sg13g2_decap_4 FILLER_50_613 ();
 sg13g2_fill_2 FILLER_50_634 ();
 sg13g2_decap_8 FILLER_50_646 ();
 sg13g2_fill_2 FILLER_50_653 ();
 sg13g2_fill_1 FILLER_50_655 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_715 ();
 sg13g2_fill_2 FILLER_50_770 ();
 sg13g2_fill_2 FILLER_50_785 ();
 sg13g2_fill_2 FILLER_50_831 ();
 sg13g2_fill_1 FILLER_50_833 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_50_892 ();
 sg13g2_decap_4 FILLER_50_918 ();
 sg13g2_fill_1 FILLER_50_922 ();
 sg13g2_decap_8 FILLER_50_930 ();
 sg13g2_decap_8 FILLER_50_941 ();
 sg13g2_decap_4 FILLER_50_948 ();
 sg13g2_fill_1 FILLER_50_978 ();
 sg13g2_fill_1 FILLER_50_1008 ();
 sg13g2_decap_4 FILLER_50_1013 ();
 sg13g2_fill_1 FILLER_50_1021 ();
 sg13g2_fill_2 FILLER_50_1041 ();
 sg13g2_fill_1 FILLER_50_1043 ();
 sg13g2_decap_8 FILLER_50_1075 ();
 sg13g2_fill_1 FILLER_50_1086 ();
 sg13g2_decap_8 FILLER_50_1091 ();
 sg13g2_fill_2 FILLER_50_1098 ();
 sg13g2_fill_1 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1110 ();
 sg13g2_decap_8 FILLER_50_1122 ();
 sg13g2_decap_8 FILLER_50_1129 ();
 sg13g2_decap_8 FILLER_50_1136 ();
 sg13g2_decap_8 FILLER_50_1143 ();
 sg13g2_decap_8 FILLER_50_1150 ();
 sg13g2_decap_8 FILLER_50_1157 ();
 sg13g2_decap_8 FILLER_50_1164 ();
 sg13g2_decap_8 FILLER_50_1171 ();
 sg13g2_decap_8 FILLER_50_1178 ();
 sg13g2_decap_8 FILLER_50_1185 ();
 sg13g2_decap_8 FILLER_50_1192 ();
 sg13g2_decap_8 FILLER_50_1199 ();
 sg13g2_decap_8 FILLER_50_1206 ();
 sg13g2_decap_8 FILLER_50_1213 ();
 sg13g2_decap_8 FILLER_50_1220 ();
 sg13g2_decap_8 FILLER_50_1227 ();
 sg13g2_decap_8 FILLER_50_1234 ();
 sg13g2_decap_8 FILLER_50_1241 ();
 sg13g2_decap_8 FILLER_50_1248 ();
 sg13g2_decap_8 FILLER_50_1255 ();
 sg13g2_decap_8 FILLER_50_1262 ();
 sg13g2_decap_8 FILLER_50_1269 ();
 sg13g2_decap_8 FILLER_50_1276 ();
 sg13g2_decap_8 FILLER_50_1283 ();
 sg13g2_decap_8 FILLER_50_1290 ();
 sg13g2_decap_8 FILLER_50_1297 ();
 sg13g2_decap_8 FILLER_50_1304 ();
 sg13g2_decap_4 FILLER_50_1311 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_4 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_60 ();
 sg13g2_decap_8 FILLER_51_88 ();
 sg13g2_decap_4 FILLER_51_95 ();
 sg13g2_fill_1 FILLER_51_99 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_4 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_149 ();
 sg13g2_fill_2 FILLER_51_178 ();
 sg13g2_decap_4 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_208 ();
 sg13g2_decap_4 FILLER_51_214 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_fill_1 FILLER_51_280 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_339 ();
 sg13g2_decap_8 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_360 ();
 sg13g2_fill_1 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_376 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_51_410 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_2 FILLER_51_475 ();
 sg13g2_fill_1 FILLER_51_477 ();
 sg13g2_fill_1 FILLER_51_492 ();
 sg13g2_decap_8 FILLER_51_510 ();
 sg13g2_fill_2 FILLER_51_517 ();
 sg13g2_fill_1 FILLER_51_519 ();
 sg13g2_fill_1 FILLER_51_524 ();
 sg13g2_fill_1 FILLER_51_551 ();
 sg13g2_fill_1 FILLER_51_557 ();
 sg13g2_decap_4 FILLER_51_562 ();
 sg13g2_fill_2 FILLER_51_566 ();
 sg13g2_fill_1 FILLER_51_580 ();
 sg13g2_decap_4 FILLER_51_589 ();
 sg13g2_fill_2 FILLER_51_593 ();
 sg13g2_decap_8 FILLER_51_599 ();
 sg13g2_fill_2 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_608 ();
 sg13g2_fill_1 FILLER_51_619 ();
 sg13g2_decap_8 FILLER_51_664 ();
 sg13g2_decap_4 FILLER_51_671 ();
 sg13g2_fill_1 FILLER_51_679 ();
 sg13g2_decap_4 FILLER_51_687 ();
 sg13g2_fill_1 FILLER_51_691 ();
 sg13g2_fill_2 FILLER_51_696 ();
 sg13g2_fill_1 FILLER_51_698 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_2 FILLER_51_736 ();
 sg13g2_decap_8 FILLER_51_743 ();
 sg13g2_decap_4 FILLER_51_750 ();
 sg13g2_decap_8 FILLER_51_802 ();
 sg13g2_decap_8 FILLER_51_809 ();
 sg13g2_fill_2 FILLER_51_816 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_fill_1 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_848 ();
 sg13g2_fill_2 FILLER_51_855 ();
 sg13g2_fill_1 FILLER_51_857 ();
 sg13g2_fill_2 FILLER_51_866 ();
 sg13g2_fill_1 FILLER_51_868 ();
 sg13g2_fill_2 FILLER_51_874 ();
 sg13g2_fill_2 FILLER_51_894 ();
 sg13g2_fill_2 FILLER_51_901 ();
 sg13g2_fill_2 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_910 ();
 sg13g2_decap_4 FILLER_51_935 ();
 sg13g2_decap_8 FILLER_51_948 ();
 sg13g2_fill_2 FILLER_51_955 ();
 sg13g2_fill_1 FILLER_51_957 ();
 sg13g2_decap_4 FILLER_51_962 ();
 sg13g2_fill_2 FILLER_51_966 ();
 sg13g2_decap_8 FILLER_51_972 ();
 sg13g2_decap_8 FILLER_51_979 ();
 sg13g2_decap_4 FILLER_51_986 ();
 sg13g2_fill_1 FILLER_51_1019 ();
 sg13g2_decap_8 FILLER_51_1038 ();
 sg13g2_fill_2 FILLER_51_1050 ();
 sg13g2_fill_2 FILLER_51_1066 ();
 sg13g2_fill_1 FILLER_51_1099 ();
 sg13g2_decap_8 FILLER_51_1126 ();
 sg13g2_decap_8 FILLER_51_1133 ();
 sg13g2_decap_8 FILLER_51_1140 ();
 sg13g2_decap_8 FILLER_51_1147 ();
 sg13g2_decap_8 FILLER_51_1154 ();
 sg13g2_decap_8 FILLER_51_1161 ();
 sg13g2_decap_8 FILLER_51_1168 ();
 sg13g2_decap_8 FILLER_51_1175 ();
 sg13g2_decap_8 FILLER_51_1182 ();
 sg13g2_decap_8 FILLER_51_1189 ();
 sg13g2_decap_8 FILLER_51_1196 ();
 sg13g2_decap_8 FILLER_51_1203 ();
 sg13g2_decap_8 FILLER_51_1210 ();
 sg13g2_decap_8 FILLER_51_1217 ();
 sg13g2_decap_8 FILLER_51_1224 ();
 sg13g2_decap_8 FILLER_51_1231 ();
 sg13g2_decap_8 FILLER_51_1238 ();
 sg13g2_decap_8 FILLER_51_1245 ();
 sg13g2_decap_8 FILLER_51_1252 ();
 sg13g2_decap_8 FILLER_51_1259 ();
 sg13g2_decap_8 FILLER_51_1266 ();
 sg13g2_decap_8 FILLER_51_1273 ();
 sg13g2_decap_8 FILLER_51_1280 ();
 sg13g2_decap_8 FILLER_51_1287 ();
 sg13g2_decap_8 FILLER_51_1294 ();
 sg13g2_decap_8 FILLER_51_1301 ();
 sg13g2_decap_8 FILLER_51_1308 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_1 FILLER_52_70 ();
 sg13g2_fill_2 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_decap_8 FILLER_52_134 ();
 sg13g2_decap_4 FILLER_52_141 ();
 sg13g2_fill_2 FILLER_52_150 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_decap_8 FILLER_52_202 ();
 sg13g2_fill_1 FILLER_52_209 ();
 sg13g2_decap_4 FILLER_52_224 ();
 sg13g2_fill_2 FILLER_52_228 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_1 FILLER_52_291 ();
 sg13g2_fill_2 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_305 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_330 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_fill_2 FILLER_52_355 ();
 sg13g2_fill_1 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_409 ();
 sg13g2_decap_4 FILLER_52_416 ();
 sg13g2_decap_4 FILLER_52_430 ();
 sg13g2_fill_1 FILLER_52_434 ();
 sg13g2_fill_1 FILLER_52_441 ();
 sg13g2_decap_4 FILLER_52_452 ();
 sg13g2_fill_1 FILLER_52_456 ();
 sg13g2_fill_2 FILLER_52_462 ();
 sg13g2_decap_4 FILLER_52_498 ();
 sg13g2_fill_2 FILLER_52_502 ();
 sg13g2_fill_2 FILLER_52_529 ();
 sg13g2_fill_1 FILLER_52_531 ();
 sg13g2_decap_4 FILLER_52_540 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_decap_4 FILLER_52_559 ();
 sg13g2_fill_2 FILLER_52_563 ();
 sg13g2_decap_4 FILLER_52_569 ();
 sg13g2_fill_2 FILLER_52_587 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_fill_1 FILLER_52_622 ();
 sg13g2_fill_2 FILLER_52_628 ();
 sg13g2_fill_1 FILLER_52_630 ();
 sg13g2_fill_2 FILLER_52_636 ();
 sg13g2_fill_1 FILLER_52_643 ();
 sg13g2_fill_2 FILLER_52_650 ();
 sg13g2_decap_4 FILLER_52_661 ();
 sg13g2_fill_1 FILLER_52_665 ();
 sg13g2_decap_4 FILLER_52_684 ();
 sg13g2_fill_2 FILLER_52_688 ();
 sg13g2_fill_2 FILLER_52_706 ();
 sg13g2_fill_2 FILLER_52_747 ();
 sg13g2_fill_1 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_755 ();
 sg13g2_fill_2 FILLER_52_762 ();
 sg13g2_fill_1 FILLER_52_764 ();
 sg13g2_fill_1 FILLER_52_769 ();
 sg13g2_decap_4 FILLER_52_850 ();
 sg13g2_decap_4 FILLER_52_919 ();
 sg13g2_fill_2 FILLER_52_923 ();
 sg13g2_fill_1 FILLER_52_951 ();
 sg13g2_fill_2 FILLER_52_983 ();
 sg13g2_fill_1 FILLER_52_985 ();
 sg13g2_decap_8 FILLER_52_990 ();
 sg13g2_decap_4 FILLER_52_997 ();
 sg13g2_fill_2 FILLER_52_1001 ();
 sg13g2_fill_1 FILLER_52_1008 ();
 sg13g2_decap_8 FILLER_52_1013 ();
 sg13g2_fill_2 FILLER_52_1020 ();
 sg13g2_fill_1 FILLER_52_1022 ();
 sg13g2_decap_4 FILLER_52_1028 ();
 sg13g2_fill_1 FILLER_52_1032 ();
 sg13g2_decap_8 FILLER_52_1037 ();
 sg13g2_decap_4 FILLER_52_1044 ();
 sg13g2_decap_4 FILLER_52_1078 ();
 sg13g2_fill_2 FILLER_52_1082 ();
 sg13g2_fill_1 FILLER_52_1088 ();
 sg13g2_decap_8 FILLER_52_1094 ();
 sg13g2_fill_2 FILLER_52_1101 ();
 sg13g2_fill_2 FILLER_52_1108 ();
 sg13g2_fill_1 FILLER_52_1110 ();
 sg13g2_decap_8 FILLER_52_1115 ();
 sg13g2_decap_8 FILLER_52_1122 ();
 sg13g2_decap_8 FILLER_52_1129 ();
 sg13g2_decap_8 FILLER_52_1136 ();
 sg13g2_decap_8 FILLER_52_1143 ();
 sg13g2_decap_8 FILLER_52_1150 ();
 sg13g2_decap_8 FILLER_52_1157 ();
 sg13g2_decap_8 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1171 ();
 sg13g2_decap_8 FILLER_52_1178 ();
 sg13g2_decap_8 FILLER_52_1185 ();
 sg13g2_decap_8 FILLER_52_1192 ();
 sg13g2_decap_8 FILLER_52_1199 ();
 sg13g2_decap_8 FILLER_52_1206 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_8 FILLER_52_1227 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_decap_8 FILLER_52_1248 ();
 sg13g2_decap_8 FILLER_52_1255 ();
 sg13g2_decap_8 FILLER_52_1262 ();
 sg13g2_decap_8 FILLER_52_1269 ();
 sg13g2_decap_8 FILLER_52_1276 ();
 sg13g2_decap_8 FILLER_52_1283 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_decap_8 FILLER_52_1297 ();
 sg13g2_decap_8 FILLER_52_1304 ();
 sg13g2_decap_4 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_71 ();
 sg13g2_decap_4 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_82 ();
 sg13g2_decap_8 FILLER_53_92 ();
 sg13g2_decap_4 FILLER_53_99 ();
 sg13g2_decap_4 FILLER_53_108 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_decap_4 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_138 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_167 ();
 sg13g2_fill_2 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_176 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_2 FILLER_53_234 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_277 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_decap_4 FILLER_53_317 ();
 sg13g2_fill_2 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_393 ();
 sg13g2_decap_4 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_decap_8 FILLER_53_440 ();
 sg13g2_fill_1 FILLER_53_447 ();
 sg13g2_decap_4 FILLER_53_482 ();
 sg13g2_decap_8 FILLER_53_491 ();
 sg13g2_fill_2 FILLER_53_498 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_fill_2 FILLER_53_525 ();
 sg13g2_decap_4 FILLER_53_553 ();
 sg13g2_fill_1 FILLER_53_583 ();
 sg13g2_fill_2 FILLER_53_606 ();
 sg13g2_fill_2 FILLER_53_612 ();
 sg13g2_fill_1 FILLER_53_629 ();
 sg13g2_fill_1 FILLER_53_637 ();
 sg13g2_fill_1 FILLER_53_648 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_decap_8 FILLER_53_662 ();
 sg13g2_decap_8 FILLER_53_669 ();
 sg13g2_fill_1 FILLER_53_676 ();
 sg13g2_decap_8 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_768 ();
 sg13g2_decap_4 FILLER_53_775 ();
 sg13g2_fill_2 FILLER_53_779 ();
 sg13g2_fill_1 FILLER_53_785 ();
 sg13g2_decap_4 FILLER_53_789 ();
 sg13g2_fill_2 FILLER_53_798 ();
 sg13g2_fill_1 FILLER_53_835 ();
 sg13g2_fill_1 FILLER_53_849 ();
 sg13g2_decap_8 FILLER_53_858 ();
 sg13g2_decap_8 FILLER_53_879 ();
 sg13g2_decap_8 FILLER_53_886 ();
 sg13g2_decap_4 FILLER_53_893 ();
 sg13g2_fill_2 FILLER_53_897 ();
 sg13g2_fill_2 FILLER_53_908 ();
 sg13g2_decap_8 FILLER_53_916 ();
 sg13g2_decap_8 FILLER_53_923 ();
 sg13g2_fill_2 FILLER_53_930 ();
 sg13g2_fill_1 FILLER_53_932 ();
 sg13g2_fill_2 FILLER_53_945 ();
 sg13g2_fill_2 FILLER_53_956 ();
 sg13g2_fill_1 FILLER_53_958 ();
 sg13g2_fill_2 FILLER_53_963 ();
 sg13g2_fill_1 FILLER_53_965 ();
 sg13g2_fill_2 FILLER_53_1053 ();
 sg13g2_decap_4 FILLER_53_1070 ();
 sg13g2_fill_1 FILLER_53_1074 ();
 sg13g2_decap_8 FILLER_53_1127 ();
 sg13g2_decap_8 FILLER_53_1134 ();
 sg13g2_decap_8 FILLER_53_1141 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1162 ();
 sg13g2_decap_8 FILLER_53_1169 ();
 sg13g2_decap_8 FILLER_53_1176 ();
 sg13g2_decap_8 FILLER_53_1183 ();
 sg13g2_decap_8 FILLER_53_1190 ();
 sg13g2_decap_8 FILLER_53_1197 ();
 sg13g2_decap_8 FILLER_53_1204 ();
 sg13g2_decap_8 FILLER_53_1211 ();
 sg13g2_decap_8 FILLER_53_1218 ();
 sg13g2_decap_8 FILLER_53_1225 ();
 sg13g2_decap_8 FILLER_53_1232 ();
 sg13g2_decap_8 FILLER_53_1239 ();
 sg13g2_decap_8 FILLER_53_1246 ();
 sg13g2_decap_8 FILLER_53_1253 ();
 sg13g2_decap_8 FILLER_53_1260 ();
 sg13g2_decap_8 FILLER_53_1267 ();
 sg13g2_decap_8 FILLER_53_1274 ();
 sg13g2_decap_8 FILLER_53_1281 ();
 sg13g2_decap_8 FILLER_53_1288 ();
 sg13g2_decap_8 FILLER_53_1295 ();
 sg13g2_decap_8 FILLER_53_1302 ();
 sg13g2_decap_4 FILLER_53_1309 ();
 sg13g2_fill_2 FILLER_53_1313 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_fill_2 FILLER_54_36 ();
 sg13g2_decap_8 FILLER_54_41 ();
 sg13g2_decap_4 FILLER_54_48 ();
 sg13g2_fill_1 FILLER_54_52 ();
 sg13g2_decap_8 FILLER_54_66 ();
 sg13g2_fill_1 FILLER_54_73 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_decap_8 FILLER_54_180 ();
 sg13g2_fill_1 FILLER_54_199 ();
 sg13g2_fill_1 FILLER_54_217 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_224 ();
 sg13g2_fill_1 FILLER_54_274 ();
 sg13g2_fill_2 FILLER_54_314 ();
 sg13g2_fill_2 FILLER_54_342 ();
 sg13g2_decap_4 FILLER_54_357 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_fill_2 FILLER_54_374 ();
 sg13g2_fill_1 FILLER_54_376 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_424 ();
 sg13g2_decap_4 FILLER_54_431 ();
 sg13g2_fill_1 FILLER_54_435 ();
 sg13g2_fill_1 FILLER_54_458 ();
 sg13g2_fill_2 FILLER_54_463 ();
 sg13g2_fill_2 FILLER_54_479 ();
 sg13g2_fill_1 FILLER_54_481 ();
 sg13g2_decap_4 FILLER_54_494 ();
 sg13g2_fill_2 FILLER_54_498 ();
 sg13g2_decap_4 FILLER_54_520 ();
 sg13g2_decap_4 FILLER_54_535 ();
 sg13g2_fill_2 FILLER_54_539 ();
 sg13g2_fill_1 FILLER_54_567 ();
 sg13g2_fill_2 FILLER_54_581 ();
 sg13g2_fill_2 FILLER_54_589 ();
 sg13g2_decap_8 FILLER_54_603 ();
 sg13g2_fill_1 FILLER_54_610 ();
 sg13g2_decap_4 FILLER_54_619 ();
 sg13g2_fill_1 FILLER_54_623 ();
 sg13g2_decap_8 FILLER_54_639 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_1 FILLER_54_695 ();
 sg13g2_fill_2 FILLER_54_709 ();
 sg13g2_fill_1 FILLER_54_711 ();
 sg13g2_fill_2 FILLER_54_725 ();
 sg13g2_fill_1 FILLER_54_727 ();
 sg13g2_fill_2 FILLER_54_748 ();
 sg13g2_fill_2 FILLER_54_754 ();
 sg13g2_fill_1 FILLER_54_756 ();
 sg13g2_fill_2 FILLER_54_777 ();
 sg13g2_fill_2 FILLER_54_802 ();
 sg13g2_fill_1 FILLER_54_804 ();
 sg13g2_fill_2 FILLER_54_829 ();
 sg13g2_decap_4 FILLER_54_860 ();
 sg13g2_fill_2 FILLER_54_895 ();
 sg13g2_fill_1 FILLER_54_902 ();
 sg13g2_fill_2 FILLER_54_910 ();
 sg13g2_fill_2 FILLER_54_916 ();
 sg13g2_decap_8 FILLER_54_996 ();
 sg13g2_decap_8 FILLER_54_1003 ();
 sg13g2_fill_2 FILLER_54_1010 ();
 sg13g2_decap_8 FILLER_54_1016 ();
 sg13g2_fill_2 FILLER_54_1023 ();
 sg13g2_fill_1 FILLER_54_1025 ();
 sg13g2_decap_4 FILLER_54_1030 ();
 sg13g2_fill_1 FILLER_54_1034 ();
 sg13g2_decap_4 FILLER_54_1065 ();
 sg13g2_decap_8 FILLER_54_1079 ();
 sg13g2_fill_2 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1092 ();
 sg13g2_decap_8 FILLER_54_1097 ();
 sg13g2_decap_8 FILLER_54_1104 ();
 sg13g2_fill_2 FILLER_54_1111 ();
 sg13g2_fill_1 FILLER_54_1113 ();
 sg13g2_decap_8 FILLER_54_1122 ();
 sg13g2_decap_8 FILLER_54_1129 ();
 sg13g2_decap_8 FILLER_54_1136 ();
 sg13g2_decap_8 FILLER_54_1143 ();
 sg13g2_decap_8 FILLER_54_1150 ();
 sg13g2_decap_8 FILLER_54_1157 ();
 sg13g2_decap_8 FILLER_54_1164 ();
 sg13g2_decap_8 FILLER_54_1171 ();
 sg13g2_decap_8 FILLER_54_1178 ();
 sg13g2_decap_8 FILLER_54_1185 ();
 sg13g2_decap_8 FILLER_54_1192 ();
 sg13g2_decap_8 FILLER_54_1199 ();
 sg13g2_decap_8 FILLER_54_1206 ();
 sg13g2_decap_8 FILLER_54_1213 ();
 sg13g2_decap_8 FILLER_54_1220 ();
 sg13g2_decap_8 FILLER_54_1227 ();
 sg13g2_decap_8 FILLER_54_1234 ();
 sg13g2_decap_8 FILLER_54_1241 ();
 sg13g2_decap_8 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1255 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_decap_8 FILLER_54_1269 ();
 sg13g2_decap_8 FILLER_54_1276 ();
 sg13g2_decap_8 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1290 ();
 sg13g2_decap_8 FILLER_54_1297 ();
 sg13g2_decap_8 FILLER_54_1304 ();
 sg13g2_decap_4 FILLER_54_1311 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_75 ();
 sg13g2_decap_4 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_117 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_fill_1 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_139 ();
 sg13g2_fill_2 FILLER_55_156 ();
 sg13g2_decap_4 FILLER_55_165 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_decap_4 FILLER_55_174 ();
 sg13g2_fill_2 FILLER_55_178 ();
 sg13g2_fill_2 FILLER_55_206 ();
 sg13g2_decap_4 FILLER_55_232 ();
 sg13g2_fill_1 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_282 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_decap_4 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_351 ();
 sg13g2_decap_4 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_55_415 ();
 sg13g2_fill_1 FILLER_55_417 ();
 sg13g2_fill_1 FILLER_55_470 ();
 sg13g2_fill_1 FILLER_55_484 ();
 sg13g2_fill_1 FILLER_55_504 ();
 sg13g2_decap_4 FILLER_55_520 ();
 sg13g2_decap_4 FILLER_55_532 ();
 sg13g2_fill_1 FILLER_55_536 ();
 sg13g2_decap_4 FILLER_55_568 ();
 sg13g2_fill_1 FILLER_55_594 ();
 sg13g2_decap_4 FILLER_55_603 ();
 sg13g2_fill_2 FILLER_55_614 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_decap_4 FILLER_55_658 ();
 sg13g2_fill_2 FILLER_55_662 ();
 sg13g2_fill_2 FILLER_55_672 ();
 sg13g2_fill_1 FILLER_55_679 ();
 sg13g2_fill_1 FILLER_55_714 ();
 sg13g2_decap_8 FILLER_55_723 ();
 sg13g2_fill_1 FILLER_55_730 ();
 sg13g2_fill_2 FILLER_55_767 ();
 sg13g2_fill_1 FILLER_55_769 ();
 sg13g2_decap_4 FILLER_55_816 ();
 sg13g2_fill_2 FILLER_55_820 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_4 FILLER_55_849 ();
 sg13g2_fill_2 FILLER_55_853 ();
 sg13g2_fill_1 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_55_866 ();
 sg13g2_decap_4 FILLER_55_881 ();
 sg13g2_fill_2 FILLER_55_931 ();
 sg13g2_decap_4 FILLER_55_945 ();
 sg13g2_decap_8 FILLER_55_957 ();
 sg13g2_decap_8 FILLER_55_969 ();
 sg13g2_decap_4 FILLER_55_976 ();
 sg13g2_fill_1 FILLER_55_980 ();
 sg13g2_decap_4 FILLER_55_985 ();
 sg13g2_fill_1 FILLER_55_989 ();
 sg13g2_fill_1 FILLER_55_1026 ();
 sg13g2_fill_1 FILLER_55_1032 ();
 sg13g2_decap_8 FILLER_55_1038 ();
 sg13g2_decap_4 FILLER_55_1054 ();
 sg13g2_fill_1 FILLER_55_1058 ();
 sg13g2_fill_2 FILLER_55_1089 ();
 sg13g2_fill_1 FILLER_55_1091 ();
 sg13g2_decap_8 FILLER_55_1116 ();
 sg13g2_decap_8 FILLER_55_1123 ();
 sg13g2_decap_8 FILLER_55_1130 ();
 sg13g2_decap_8 FILLER_55_1137 ();
 sg13g2_decap_8 FILLER_55_1144 ();
 sg13g2_decap_8 FILLER_55_1151 ();
 sg13g2_decap_8 FILLER_55_1158 ();
 sg13g2_decap_8 FILLER_55_1165 ();
 sg13g2_decap_8 FILLER_55_1172 ();
 sg13g2_decap_8 FILLER_55_1179 ();
 sg13g2_decap_8 FILLER_55_1186 ();
 sg13g2_decap_8 FILLER_55_1193 ();
 sg13g2_decap_8 FILLER_55_1200 ();
 sg13g2_decap_8 FILLER_55_1207 ();
 sg13g2_decap_8 FILLER_55_1214 ();
 sg13g2_decap_8 FILLER_55_1221 ();
 sg13g2_decap_8 FILLER_55_1228 ();
 sg13g2_decap_8 FILLER_55_1235 ();
 sg13g2_decap_8 FILLER_55_1242 ();
 sg13g2_decap_8 FILLER_55_1249 ();
 sg13g2_decap_8 FILLER_55_1256 ();
 sg13g2_decap_8 FILLER_55_1263 ();
 sg13g2_decap_8 FILLER_55_1270 ();
 sg13g2_decap_8 FILLER_55_1277 ();
 sg13g2_decap_8 FILLER_55_1284 ();
 sg13g2_decap_8 FILLER_55_1291 ();
 sg13g2_decap_8 FILLER_55_1298 ();
 sg13g2_decap_8 FILLER_55_1305 ();
 sg13g2_fill_2 FILLER_55_1312 ();
 sg13g2_fill_1 FILLER_55_1314 ();
 sg13g2_fill_2 FILLER_56_26 ();
 sg13g2_decap_8 FILLER_56_50 ();
 sg13g2_decap_4 FILLER_56_57 ();
 sg13g2_fill_1 FILLER_56_61 ();
 sg13g2_decap_8 FILLER_56_107 ();
 sg13g2_fill_1 FILLER_56_114 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_185 ();
 sg13g2_decap_8 FILLER_56_190 ();
 sg13g2_fill_2 FILLER_56_197 ();
 sg13g2_decap_4 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_208 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_296 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_fill_1 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_349 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_decap_4 FILLER_56_357 ();
 sg13g2_decap_4 FILLER_56_365 ();
 sg13g2_decap_4 FILLER_56_373 ();
 sg13g2_decap_4 FILLER_56_414 ();
 sg13g2_decap_8 FILLER_56_440 ();
 sg13g2_decap_4 FILLER_56_447 ();
 sg13g2_decap_8 FILLER_56_470 ();
 sg13g2_fill_2 FILLER_56_477 ();
 sg13g2_decap_4 FILLER_56_487 ();
 sg13g2_fill_1 FILLER_56_491 ();
 sg13g2_fill_2 FILLER_56_508 ();
 sg13g2_decap_8 FILLER_56_515 ();
 sg13g2_fill_1 FILLER_56_522 ();
 sg13g2_decap_8 FILLER_56_533 ();
 sg13g2_fill_1 FILLER_56_545 ();
 sg13g2_fill_2 FILLER_56_559 ();
 sg13g2_fill_1 FILLER_56_561 ();
 sg13g2_decap_4 FILLER_56_578 ();
 sg13g2_fill_2 FILLER_56_592 ();
 sg13g2_decap_8 FILLER_56_599 ();
 sg13g2_fill_2 FILLER_56_606 ();
 sg13g2_fill_1 FILLER_56_608 ();
 sg13g2_fill_2 FILLER_56_617 ();
 sg13g2_fill_1 FILLER_56_619 ();
 sg13g2_fill_1 FILLER_56_632 ();
 sg13g2_fill_1 FILLER_56_656 ();
 sg13g2_decap_8 FILLER_56_672 ();
 sg13g2_fill_2 FILLER_56_687 ();
 sg13g2_fill_1 FILLER_56_725 ();
 sg13g2_decap_8 FILLER_56_740 ();
 sg13g2_decap_4 FILLER_56_747 ();
 sg13g2_fill_1 FILLER_56_751 ();
 sg13g2_decap_4 FILLER_56_756 ();
 sg13g2_fill_1 FILLER_56_770 ();
 sg13g2_decap_4 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_798 ();
 sg13g2_decap_4 FILLER_56_814 ();
 sg13g2_fill_1 FILLER_56_818 ();
 sg13g2_fill_2 FILLER_56_829 ();
 sg13g2_decap_4 FILLER_56_867 ();
 sg13g2_fill_2 FILLER_56_925 ();
 sg13g2_fill_2 FILLER_56_953 ();
 sg13g2_fill_2 FILLER_56_991 ();
 sg13g2_fill_1 FILLER_56_993 ();
 sg13g2_decap_8 FILLER_56_1019 ();
 sg13g2_fill_1 FILLER_56_1042 ();
 sg13g2_decap_4 FILLER_56_1048 ();
 sg13g2_decap_4 FILLER_56_1063 ();
 sg13g2_fill_1 FILLER_56_1067 ();
 sg13g2_decap_8 FILLER_56_1113 ();
 sg13g2_decap_8 FILLER_56_1120 ();
 sg13g2_decap_8 FILLER_56_1127 ();
 sg13g2_decap_8 FILLER_56_1134 ();
 sg13g2_decap_8 FILLER_56_1141 ();
 sg13g2_decap_8 FILLER_56_1148 ();
 sg13g2_decap_8 FILLER_56_1155 ();
 sg13g2_decap_8 FILLER_56_1162 ();
 sg13g2_decap_8 FILLER_56_1169 ();
 sg13g2_decap_8 FILLER_56_1176 ();
 sg13g2_decap_8 FILLER_56_1183 ();
 sg13g2_decap_8 FILLER_56_1190 ();
 sg13g2_decap_8 FILLER_56_1197 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1218 ();
 sg13g2_decap_8 FILLER_56_1225 ();
 sg13g2_decap_8 FILLER_56_1232 ();
 sg13g2_decap_8 FILLER_56_1239 ();
 sg13g2_decap_8 FILLER_56_1246 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1267 ();
 sg13g2_decap_8 FILLER_56_1274 ();
 sg13g2_decap_8 FILLER_56_1281 ();
 sg13g2_decap_8 FILLER_56_1288 ();
 sg13g2_decap_8 FILLER_56_1295 ();
 sg13g2_decap_8 FILLER_56_1302 ();
 sg13g2_decap_4 FILLER_56_1309 ();
 sg13g2_fill_2 FILLER_56_1313 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_18 ();
 sg13g2_decap_8 FILLER_57_43 ();
 sg13g2_decap_4 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_54 ();
 sg13g2_decap_8 FILLER_57_65 ();
 sg13g2_decap_8 FILLER_57_72 ();
 sg13g2_decap_8 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_125 ();
 sg13g2_decap_4 FILLER_57_132 ();
 sg13g2_decap_8 FILLER_57_145 ();
 sg13g2_fill_2 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_167 ();
 sg13g2_decap_8 FILLER_57_174 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_fill_2 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_2 FILLER_57_278 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_fill_2 FILLER_57_313 ();
 sg13g2_fill_1 FILLER_57_331 ();
 sg13g2_decap_4 FILLER_57_356 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_fill_1 FILLER_57_417 ();
 sg13g2_fill_2 FILLER_57_423 ();
 sg13g2_decap_8 FILLER_57_451 ();
 sg13g2_decap_4 FILLER_57_458 ();
 sg13g2_fill_1 FILLER_57_462 ();
 sg13g2_fill_2 FILLER_57_479 ();
 sg13g2_fill_1 FILLER_57_481 ();
 sg13g2_decap_8 FILLER_57_485 ();
 sg13g2_decap_8 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_499 ();
 sg13g2_fill_2 FILLER_57_504 ();
 sg13g2_decap_4 FILLER_57_514 ();
 sg13g2_decap_4 FILLER_57_544 ();
 sg13g2_decap_4 FILLER_57_555 ();
 sg13g2_fill_2 FILLER_57_559 ();
 sg13g2_fill_2 FILLER_57_578 ();
 sg13g2_fill_1 FILLER_57_580 ();
 sg13g2_decap_8 FILLER_57_601 ();
 sg13g2_decap_4 FILLER_57_608 ();
 sg13g2_fill_2 FILLER_57_612 ();
 sg13g2_decap_8 FILLER_57_618 ();
 sg13g2_fill_1 FILLER_57_625 ();
 sg13g2_fill_1 FILLER_57_631 ();
 sg13g2_decap_8 FILLER_57_638 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_decap_8 FILLER_57_650 ();
 sg13g2_fill_1 FILLER_57_657 ();
 sg13g2_fill_2 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_decap_8 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_703 ();
 sg13g2_fill_2 FILLER_57_710 ();
 sg13g2_fill_1 FILLER_57_712 ();
 sg13g2_fill_1 FILLER_57_722 ();
 sg13g2_fill_2 FILLER_57_785 ();
 sg13g2_decap_8 FILLER_57_813 ();
 sg13g2_fill_2 FILLER_57_820 ();
 sg13g2_fill_2 FILLER_57_848 ();
 sg13g2_fill_1 FILLER_57_850 ();
 sg13g2_fill_2 FILLER_57_855 ();
 sg13g2_fill_1 FILLER_57_864 ();
 sg13g2_decap_8 FILLER_57_873 ();
 sg13g2_fill_2 FILLER_57_880 ();
 sg13g2_fill_2 FILLER_57_886 ();
 sg13g2_fill_1 FILLER_57_906 ();
 sg13g2_decap_4 FILLER_57_933 ();
 sg13g2_fill_1 FILLER_57_937 ();
 sg13g2_fill_2 FILLER_57_942 ();
 sg13g2_fill_2 FILLER_57_959 ();
 sg13g2_fill_2 FILLER_57_1031 ();
 sg13g2_fill_1 FILLER_57_1033 ();
 sg13g2_fill_2 FILLER_57_1052 ();
 sg13g2_fill_1 FILLER_57_1105 ();
 sg13g2_decap_8 FILLER_57_1110 ();
 sg13g2_decap_8 FILLER_57_1117 ();
 sg13g2_decap_8 FILLER_57_1124 ();
 sg13g2_decap_8 FILLER_57_1131 ();
 sg13g2_decap_8 FILLER_57_1138 ();
 sg13g2_decap_8 FILLER_57_1145 ();
 sg13g2_decap_8 FILLER_57_1152 ();
 sg13g2_decap_8 FILLER_57_1159 ();
 sg13g2_decap_8 FILLER_57_1166 ();
 sg13g2_decap_8 FILLER_57_1173 ();
 sg13g2_decap_8 FILLER_57_1180 ();
 sg13g2_decap_8 FILLER_57_1187 ();
 sg13g2_decap_8 FILLER_57_1194 ();
 sg13g2_decap_8 FILLER_57_1201 ();
 sg13g2_decap_8 FILLER_57_1208 ();
 sg13g2_decap_8 FILLER_57_1215 ();
 sg13g2_decap_8 FILLER_57_1222 ();
 sg13g2_decap_8 FILLER_57_1229 ();
 sg13g2_decap_8 FILLER_57_1236 ();
 sg13g2_decap_8 FILLER_57_1243 ();
 sg13g2_decap_8 FILLER_57_1250 ();
 sg13g2_decap_8 FILLER_57_1257 ();
 sg13g2_decap_8 FILLER_57_1264 ();
 sg13g2_decap_8 FILLER_57_1271 ();
 sg13g2_decap_8 FILLER_57_1278 ();
 sg13g2_decap_8 FILLER_57_1285 ();
 sg13g2_decap_8 FILLER_57_1292 ();
 sg13g2_decap_8 FILLER_57_1299 ();
 sg13g2_decap_8 FILLER_57_1306 ();
 sg13g2_fill_2 FILLER_57_1313 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_27 ();
 sg13g2_fill_1 FILLER_58_31 ();
 sg13g2_decap_4 FILLER_58_39 ();
 sg13g2_fill_2 FILLER_58_43 ();
 sg13g2_fill_1 FILLER_58_57 ();
 sg13g2_fill_1 FILLER_58_95 ();
 sg13g2_decap_4 FILLER_58_127 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_192 ();
 sg13g2_decap_4 FILLER_58_212 ();
 sg13g2_decap_4 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_308 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_decap_4 FILLER_58_337 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_decap_4 FILLER_58_358 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_2 FILLER_58_371 ();
 sg13g2_fill_1 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_424 ();
 sg13g2_fill_2 FILLER_58_460 ();
 sg13g2_fill_2 FILLER_58_472 ();
 sg13g2_decap_8 FILLER_58_514 ();
 sg13g2_fill_2 FILLER_58_521 ();
 sg13g2_fill_1 FILLER_58_537 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_decap_4 FILLER_58_567 ();
 sg13g2_fill_2 FILLER_58_601 ();
 sg13g2_fill_2 FILLER_58_629 ();
 sg13g2_decap_8 FILLER_58_657 ();
 sg13g2_decap_8 FILLER_58_664 ();
 sg13g2_decap_4 FILLER_58_679 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_fill_1 FILLER_58_711 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_748 ();
 sg13g2_decap_8 FILLER_58_753 ();
 sg13g2_decap_8 FILLER_58_760 ();
 sg13g2_decap_8 FILLER_58_767 ();
 sg13g2_decap_8 FILLER_58_774 ();
 sg13g2_decap_8 FILLER_58_781 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_fill_2 FILLER_58_795 ();
 sg13g2_fill_1 FILLER_58_797 ();
 sg13g2_decap_8 FILLER_58_810 ();
 sg13g2_decap_4 FILLER_58_817 ();
 sg13g2_fill_1 FILLER_58_831 ();
 sg13g2_decap_8 FILLER_58_836 ();
 sg13g2_decap_4 FILLER_58_843 ();
 sg13g2_fill_1 FILLER_58_859 ();
 sg13g2_fill_2 FILLER_58_865 ();
 sg13g2_decap_8 FILLER_58_882 ();
 sg13g2_decap_8 FILLER_58_904 ();
 sg13g2_decap_8 FILLER_58_911 ();
 sg13g2_decap_4 FILLER_58_922 ();
 sg13g2_fill_2 FILLER_58_926 ();
 sg13g2_decap_8 FILLER_58_937 ();
 sg13g2_fill_2 FILLER_58_944 ();
 sg13g2_fill_1 FILLER_58_960 ();
 sg13g2_decap_8 FILLER_58_969 ();
 sg13g2_fill_2 FILLER_58_980 ();
 sg13g2_decap_8 FILLER_58_986 ();
 sg13g2_decap_8 FILLER_58_993 ();
 sg13g2_decap_4 FILLER_58_1000 ();
 sg13g2_fill_2 FILLER_58_1004 ();
 sg13g2_fill_2 FILLER_58_1015 ();
 sg13g2_fill_1 FILLER_58_1017 ();
 sg13g2_fill_1 FILLER_58_1041 ();
 sg13g2_fill_2 FILLER_58_1047 ();
 sg13g2_decap_8 FILLER_58_1064 ();
 sg13g2_decap_8 FILLER_58_1071 ();
 sg13g2_fill_2 FILLER_58_1078 ();
 sg13g2_decap_8 FILLER_58_1084 ();
 sg13g2_decap_4 FILLER_58_1091 ();
 sg13g2_decap_8 FILLER_58_1121 ();
 sg13g2_decap_8 FILLER_58_1128 ();
 sg13g2_decap_8 FILLER_58_1135 ();
 sg13g2_decap_8 FILLER_58_1142 ();
 sg13g2_decap_8 FILLER_58_1149 ();
 sg13g2_decap_8 FILLER_58_1156 ();
 sg13g2_decap_8 FILLER_58_1163 ();
 sg13g2_decap_8 FILLER_58_1170 ();
 sg13g2_decap_8 FILLER_58_1177 ();
 sg13g2_decap_8 FILLER_58_1184 ();
 sg13g2_decap_8 FILLER_58_1191 ();
 sg13g2_decap_8 FILLER_58_1198 ();
 sg13g2_decap_8 FILLER_58_1205 ();
 sg13g2_decap_8 FILLER_58_1212 ();
 sg13g2_decap_8 FILLER_58_1219 ();
 sg13g2_decap_8 FILLER_58_1226 ();
 sg13g2_decap_8 FILLER_58_1233 ();
 sg13g2_decap_8 FILLER_58_1240 ();
 sg13g2_decap_8 FILLER_58_1247 ();
 sg13g2_decap_8 FILLER_58_1254 ();
 sg13g2_decap_8 FILLER_58_1261 ();
 sg13g2_decap_8 FILLER_58_1268 ();
 sg13g2_decap_8 FILLER_58_1275 ();
 sg13g2_decap_8 FILLER_58_1282 ();
 sg13g2_decap_8 FILLER_58_1289 ();
 sg13g2_decap_8 FILLER_58_1296 ();
 sg13g2_decap_8 FILLER_58_1303 ();
 sg13g2_decap_4 FILLER_58_1310 ();
 sg13g2_fill_1 FILLER_58_1314 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_4 ();
 sg13g2_decap_4 FILLER_59_9 ();
 sg13g2_decap_8 FILLER_59_71 ();
 sg13g2_decap_4 FILLER_59_78 ();
 sg13g2_fill_1 FILLER_59_82 ();
 sg13g2_fill_2 FILLER_59_101 ();
 sg13g2_decap_4 FILLER_59_109 ();
 sg13g2_decap_8 FILLER_59_122 ();
 sg13g2_decap_4 FILLER_59_137 ();
 sg13g2_fill_2 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_4 FILLER_59_179 ();
 sg13g2_fill_2 FILLER_59_183 ();
 sg13g2_decap_4 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_237 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_312 ();
 sg13g2_fill_1 FILLER_59_314 ();
 sg13g2_fill_1 FILLER_59_337 ();
 sg13g2_decap_8 FILLER_59_344 ();
 sg13g2_decap_4 FILLER_59_351 ();
 sg13g2_fill_2 FILLER_59_355 ();
 sg13g2_fill_2 FILLER_59_371 ();
 sg13g2_fill_2 FILLER_59_377 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_fill_1 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_fill_1 FILLER_59_435 ();
 sg13g2_decap_8 FILLER_59_443 ();
 sg13g2_decap_4 FILLER_59_466 ();
 sg13g2_fill_2 FILLER_59_475 ();
 sg13g2_fill_2 FILLER_59_487 ();
 sg13g2_fill_1 FILLER_59_489 ();
 sg13g2_fill_1 FILLER_59_494 ();
 sg13g2_fill_1 FILLER_59_509 ();
 sg13g2_decap_8 FILLER_59_536 ();
 sg13g2_decap_4 FILLER_59_543 ();
 sg13g2_fill_1 FILLER_59_547 ();
 sg13g2_fill_1 FILLER_59_586 ();
 sg13g2_fill_2 FILLER_59_597 ();
 sg13g2_decap_4 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_639 ();
 sg13g2_fill_2 FILLER_59_692 ();
 sg13g2_decap_8 FILLER_59_698 ();
 sg13g2_decap_8 FILLER_59_705 ();
 sg13g2_fill_2 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_771 ();
 sg13g2_fill_1 FILLER_59_777 ();
 sg13g2_fill_1 FILLER_59_787 ();
 sg13g2_decap_8 FILLER_59_793 ();
 sg13g2_fill_1 FILLER_59_805 ();
 sg13g2_fill_2 FILLER_59_811 ();
 sg13g2_fill_2 FILLER_59_867 ();
 sg13g2_decap_8 FILLER_59_913 ();
 sg13g2_fill_2 FILLER_59_920 ();
 sg13g2_fill_2 FILLER_59_935 ();
 sg13g2_fill_2 FILLER_59_1023 ();
 sg13g2_fill_1 FILLER_59_1025 ();
 sg13g2_fill_2 FILLER_59_1035 ();
 sg13g2_fill_2 FILLER_59_1061 ();
 sg13g2_decap_4 FILLER_59_1099 ();
 sg13g2_fill_2 FILLER_59_1103 ();
 sg13g2_fill_1 FILLER_59_1109 ();
 sg13g2_decap_8 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1120 ();
 sg13g2_decap_8 FILLER_59_1127 ();
 sg13g2_decap_8 FILLER_59_1134 ();
 sg13g2_decap_8 FILLER_59_1141 ();
 sg13g2_decap_8 FILLER_59_1148 ();
 sg13g2_decap_8 FILLER_59_1155 ();
 sg13g2_decap_8 FILLER_59_1162 ();
 sg13g2_decap_8 FILLER_59_1169 ();
 sg13g2_decap_8 FILLER_59_1176 ();
 sg13g2_decap_8 FILLER_59_1183 ();
 sg13g2_decap_8 FILLER_59_1190 ();
 sg13g2_decap_8 FILLER_59_1197 ();
 sg13g2_decap_8 FILLER_59_1204 ();
 sg13g2_decap_8 FILLER_59_1211 ();
 sg13g2_decap_8 FILLER_59_1218 ();
 sg13g2_decap_8 FILLER_59_1225 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_8 FILLER_59_1253 ();
 sg13g2_decap_8 FILLER_59_1260 ();
 sg13g2_decap_8 FILLER_59_1267 ();
 sg13g2_decap_8 FILLER_59_1274 ();
 sg13g2_decap_8 FILLER_59_1281 ();
 sg13g2_decap_8 FILLER_59_1288 ();
 sg13g2_decap_8 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1302 ();
 sg13g2_decap_4 FILLER_59_1309 ();
 sg13g2_fill_2 FILLER_59_1313 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_60 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_167 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_211 ();
 sg13g2_decap_8 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_244 ();
 sg13g2_decap_8 FILLER_60_262 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_324 ();
 sg13g2_decap_4 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_412 ();
 sg13g2_fill_1 FILLER_60_439 ();
 sg13g2_decap_4 FILLER_60_456 ();
 sg13g2_fill_1 FILLER_60_460 ();
 sg13g2_decap_4 FILLER_60_472 ();
 sg13g2_fill_1 FILLER_60_476 ();
 sg13g2_decap_4 FILLER_60_486 ();
 sg13g2_fill_2 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_496 ();
 sg13g2_fill_2 FILLER_60_506 ();
 sg13g2_fill_1 FILLER_60_508 ();
 sg13g2_fill_1 FILLER_60_519 ();
 sg13g2_decap_8 FILLER_60_524 ();
 sg13g2_decap_4 FILLER_60_531 ();
 sg13g2_decap_4 FILLER_60_539 ();
 sg13g2_decap_8 FILLER_60_568 ();
 sg13g2_decap_4 FILLER_60_587 ();
 sg13g2_fill_2 FILLER_60_591 ();
 sg13g2_fill_2 FILLER_60_616 ();
 sg13g2_fill_1 FILLER_60_618 ();
 sg13g2_fill_2 FILLER_60_627 ();
 sg13g2_fill_1 FILLER_60_629 ();
 sg13g2_fill_1 FILLER_60_634 ();
 sg13g2_decap_4 FILLER_60_662 ();
 sg13g2_fill_2 FILLER_60_674 ();
 sg13g2_fill_1 FILLER_60_680 ();
 sg13g2_decap_8 FILLER_60_726 ();
 sg13g2_decap_8 FILLER_60_733 ();
 sg13g2_fill_2 FILLER_60_748 ();
 sg13g2_decap_8 FILLER_60_772 ();
 sg13g2_decap_4 FILLER_60_779 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_8 FILLER_60_820 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_fill_1 FILLER_60_852 ();
 sg13g2_decap_8 FILLER_60_866 ();
 sg13g2_decap_4 FILLER_60_873 ();
 sg13g2_fill_2 FILLER_60_877 ();
 sg13g2_decap_4 FILLER_60_883 ();
 sg13g2_fill_2 FILLER_60_893 ();
 sg13g2_fill_2 FILLER_60_912 ();
 sg13g2_fill_1 FILLER_60_914 ();
 sg13g2_fill_2 FILLER_60_944 ();
 sg13g2_fill_2 FILLER_60_963 ();
 sg13g2_decap_8 FILLER_60_975 ();
 sg13g2_fill_1 FILLER_60_982 ();
 sg13g2_fill_2 FILLER_60_987 ();
 sg13g2_decap_4 FILLER_60_999 ();
 sg13g2_fill_1 FILLER_60_1003 ();
 sg13g2_decap_4 FILLER_60_1008 ();
 sg13g2_decap_8 FILLER_60_1022 ();
 sg13g2_decap_4 FILLER_60_1038 ();
 sg13g2_fill_2 FILLER_60_1042 ();
 sg13g2_fill_2 FILLER_60_1049 ();
 sg13g2_decap_8 FILLER_60_1061 ();
 sg13g2_fill_1 FILLER_60_1068 ();
 sg13g2_fill_2 FILLER_60_1072 ();
 sg13g2_fill_2 FILLER_60_1081 ();
 sg13g2_fill_1 FILLER_60_1083 ();
 sg13g2_decap_8 FILLER_60_1120 ();
 sg13g2_decap_8 FILLER_60_1127 ();
 sg13g2_decap_8 FILLER_60_1134 ();
 sg13g2_decap_8 FILLER_60_1141 ();
 sg13g2_decap_8 FILLER_60_1148 ();
 sg13g2_decap_8 FILLER_60_1155 ();
 sg13g2_decap_8 FILLER_60_1162 ();
 sg13g2_decap_8 FILLER_60_1169 ();
 sg13g2_decap_8 FILLER_60_1176 ();
 sg13g2_decap_8 FILLER_60_1183 ();
 sg13g2_decap_8 FILLER_60_1190 ();
 sg13g2_decap_8 FILLER_60_1197 ();
 sg13g2_decap_8 FILLER_60_1204 ();
 sg13g2_decap_8 FILLER_60_1211 ();
 sg13g2_decap_8 FILLER_60_1218 ();
 sg13g2_decap_8 FILLER_60_1225 ();
 sg13g2_decap_8 FILLER_60_1232 ();
 sg13g2_decap_8 FILLER_60_1239 ();
 sg13g2_decap_8 FILLER_60_1246 ();
 sg13g2_decap_8 FILLER_60_1253 ();
 sg13g2_decap_8 FILLER_60_1260 ();
 sg13g2_decap_8 FILLER_60_1267 ();
 sg13g2_decap_8 FILLER_60_1274 ();
 sg13g2_decap_8 FILLER_60_1281 ();
 sg13g2_decap_8 FILLER_60_1288 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_8 FILLER_60_1302 ();
 sg13g2_decap_4 FILLER_60_1309 ();
 sg13g2_fill_2 FILLER_60_1313 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_4 ();
 sg13g2_fill_1 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_19 ();
 sg13g2_fill_2 FILLER_61_26 ();
 sg13g2_fill_1 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_41 ();
 sg13g2_decap_8 FILLER_61_51 ();
 sg13g2_decap_8 FILLER_61_58 ();
 sg13g2_decap_4 FILLER_61_65 ();
 sg13g2_fill_2 FILLER_61_100 ();
 sg13g2_fill_1 FILLER_61_102 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_fill_1 FILLER_61_136 ();
 sg13g2_decap_4 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_144 ();
 sg13g2_fill_1 FILLER_61_150 ();
 sg13g2_decap_8 FILLER_61_155 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_170 ();
 sg13g2_decap_4 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_fill_2 FILLER_61_228 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_fill_2 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_352 ();
 sg13g2_decap_8 FILLER_61_366 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_380 ();
 sg13g2_fill_2 FILLER_61_386 ();
 sg13g2_decap_4 FILLER_61_414 ();
 sg13g2_fill_1 FILLER_61_418 ();
 sg13g2_decap_8 FILLER_61_423 ();
 sg13g2_fill_1 FILLER_61_430 ();
 sg13g2_decap_8 FILLER_61_440 ();
 sg13g2_fill_1 FILLER_61_447 ();
 sg13g2_fill_1 FILLER_61_453 ();
 sg13g2_decap_4 FILLER_61_475 ();
 sg13g2_decap_4 FILLER_61_521 ();
 sg13g2_decap_4 FILLER_61_551 ();
 sg13g2_decap_8 FILLER_61_565 ();
 sg13g2_fill_2 FILLER_61_572 ();
 sg13g2_decap_4 FILLER_61_579 ();
 sg13g2_decap_4 FILLER_61_614 ();
 sg13g2_fill_1 FILLER_61_618 ();
 sg13g2_decap_8 FILLER_61_645 ();
 sg13g2_fill_1 FILLER_61_656 ();
 sg13g2_decap_8 FILLER_61_661 ();
 sg13g2_fill_2 FILLER_61_668 ();
 sg13g2_decap_4 FILLER_61_706 ();
 sg13g2_fill_1 FILLER_61_710 ();
 sg13g2_fill_1 FILLER_61_715 ();
 sg13g2_decap_8 FILLER_61_720 ();
 sg13g2_fill_2 FILLER_61_727 ();
 sg13g2_fill_1 FILLER_61_729 ();
 sg13g2_decap_4 FILLER_61_740 ();
 sg13g2_fill_2 FILLER_61_744 ();
 sg13g2_fill_2 FILLER_61_760 ();
 sg13g2_decap_8 FILLER_61_798 ();
 sg13g2_decap_4 FILLER_61_809 ();
 sg13g2_fill_1 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_854 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_61_898 ();
 sg13g2_decap_8 FILLER_61_905 ();
 sg13g2_decap_8 FILLER_61_912 ();
 sg13g2_fill_2 FILLER_61_919 ();
 sg13g2_fill_1 FILLER_61_921 ();
 sg13g2_fill_1 FILLER_61_937 ();
 sg13g2_decap_8 FILLER_61_964 ();
 sg13g2_fill_2 FILLER_61_1090 ();
 sg13g2_decap_8 FILLER_61_1121 ();
 sg13g2_decap_8 FILLER_61_1128 ();
 sg13g2_decap_8 FILLER_61_1135 ();
 sg13g2_decap_8 FILLER_61_1142 ();
 sg13g2_decap_8 FILLER_61_1149 ();
 sg13g2_decap_8 FILLER_61_1156 ();
 sg13g2_decap_8 FILLER_61_1163 ();
 sg13g2_decap_8 FILLER_61_1170 ();
 sg13g2_decap_8 FILLER_61_1177 ();
 sg13g2_decap_8 FILLER_61_1184 ();
 sg13g2_decap_8 FILLER_61_1191 ();
 sg13g2_decap_8 FILLER_61_1198 ();
 sg13g2_decap_8 FILLER_61_1205 ();
 sg13g2_decap_8 FILLER_61_1212 ();
 sg13g2_decap_8 FILLER_61_1219 ();
 sg13g2_decap_8 FILLER_61_1226 ();
 sg13g2_decap_8 FILLER_61_1233 ();
 sg13g2_decap_8 FILLER_61_1240 ();
 sg13g2_decap_8 FILLER_61_1247 ();
 sg13g2_decap_8 FILLER_61_1254 ();
 sg13g2_decap_8 FILLER_61_1261 ();
 sg13g2_decap_8 FILLER_61_1268 ();
 sg13g2_decap_8 FILLER_61_1275 ();
 sg13g2_decap_8 FILLER_61_1282 ();
 sg13g2_decap_8 FILLER_61_1289 ();
 sg13g2_decap_8 FILLER_61_1296 ();
 sg13g2_decap_8 FILLER_61_1303 ();
 sg13g2_decap_4 FILLER_61_1310 ();
 sg13g2_fill_1 FILLER_61_1314 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_71 ();
 sg13g2_fill_2 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_fill_2 FILLER_62_85 ();
 sg13g2_decap_4 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_decap_8 FILLER_62_114 ();
 sg13g2_decap_8 FILLER_62_121 ();
 sg13g2_fill_2 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_156 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_2 FILLER_62_226 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_decap_4 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_317 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_325 ();
 sg13g2_fill_2 FILLER_62_369 ();
 sg13g2_fill_1 FILLER_62_378 ();
 sg13g2_fill_2 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_62_414 ();
 sg13g2_fill_2 FILLER_62_421 ();
 sg13g2_fill_1 FILLER_62_423 ();
 sg13g2_fill_1 FILLER_62_451 ();
 sg13g2_fill_1 FILLER_62_468 ();
 sg13g2_fill_1 FILLER_62_474 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_fill_2 FILLER_62_500 ();
 sg13g2_fill_1 FILLER_62_502 ();
 sg13g2_fill_2 FILLER_62_546 ();
 sg13g2_fill_1 FILLER_62_548 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_fill_1 FILLER_62_556 ();
 sg13g2_fill_2 FILLER_62_561 ();
 sg13g2_fill_1 FILLER_62_563 ();
 sg13g2_decap_8 FILLER_62_587 ();
 sg13g2_decap_4 FILLER_62_594 ();
 sg13g2_fill_1 FILLER_62_598 ();
 sg13g2_decap_8 FILLER_62_603 ();
 sg13g2_decap_4 FILLER_62_610 ();
 sg13g2_fill_2 FILLER_62_614 ();
 sg13g2_decap_4 FILLER_62_624 ();
 sg13g2_decap_4 FILLER_62_642 ();
 sg13g2_fill_1 FILLER_62_694 ();
 sg13g2_fill_2 FILLER_62_731 ();
 sg13g2_decap_8 FILLER_62_764 ();
 sg13g2_decap_8 FILLER_62_771 ();
 sg13g2_fill_2 FILLER_62_829 ();
 sg13g2_fill_1 FILLER_62_839 ();
 sg13g2_fill_2 FILLER_62_879 ();
 sg13g2_fill_1 FILLER_62_881 ();
 sg13g2_decap_8 FILLER_62_886 ();
 sg13g2_fill_1 FILLER_62_893 ();
 sg13g2_decap_8 FILLER_62_902 ();
 sg13g2_decap_4 FILLER_62_909 ();
 sg13g2_fill_1 FILLER_62_913 ();
 sg13g2_decap_4 FILLER_62_941 ();
 sg13g2_fill_1 FILLER_62_945 ();
 sg13g2_fill_1 FILLER_62_951 ();
 sg13g2_decap_4 FILLER_62_957 ();
 sg13g2_fill_1 FILLER_62_961 ();
 sg13g2_fill_1 FILLER_62_967 ();
 sg13g2_decap_8 FILLER_62_972 ();
 sg13g2_fill_2 FILLER_62_979 ();
 sg13g2_fill_1 FILLER_62_981 ();
 sg13g2_decap_8 FILLER_62_986 ();
 sg13g2_decap_4 FILLER_62_997 ();
 sg13g2_fill_2 FILLER_62_1001 ();
 sg13g2_decap_8 FILLER_62_1012 ();
 sg13g2_decap_8 FILLER_62_1019 ();
 sg13g2_decap_4 FILLER_62_1026 ();
 sg13g2_fill_1 FILLER_62_1030 ();
 sg13g2_decap_4 FILLER_62_1046 ();
 sg13g2_fill_2 FILLER_62_1055 ();
 sg13g2_fill_1 FILLER_62_1057 ();
 sg13g2_decap_8 FILLER_62_1072 ();
 sg13g2_decap_8 FILLER_62_1079 ();
 sg13g2_decap_8 FILLER_62_1096 ();
 sg13g2_decap_8 FILLER_62_1107 ();
 sg13g2_decap_8 FILLER_62_1114 ();
 sg13g2_decap_8 FILLER_62_1121 ();
 sg13g2_decap_8 FILLER_62_1128 ();
 sg13g2_decap_8 FILLER_62_1135 ();
 sg13g2_decap_8 FILLER_62_1142 ();
 sg13g2_decap_8 FILLER_62_1149 ();
 sg13g2_decap_8 FILLER_62_1156 ();
 sg13g2_decap_8 FILLER_62_1163 ();
 sg13g2_decap_8 FILLER_62_1170 ();
 sg13g2_decap_8 FILLER_62_1177 ();
 sg13g2_decap_8 FILLER_62_1184 ();
 sg13g2_decap_8 FILLER_62_1191 ();
 sg13g2_decap_8 FILLER_62_1198 ();
 sg13g2_decap_8 FILLER_62_1205 ();
 sg13g2_decap_8 FILLER_62_1212 ();
 sg13g2_decap_8 FILLER_62_1219 ();
 sg13g2_decap_8 FILLER_62_1226 ();
 sg13g2_decap_8 FILLER_62_1233 ();
 sg13g2_decap_8 FILLER_62_1240 ();
 sg13g2_decap_8 FILLER_62_1247 ();
 sg13g2_decap_8 FILLER_62_1254 ();
 sg13g2_decap_8 FILLER_62_1261 ();
 sg13g2_decap_8 FILLER_62_1268 ();
 sg13g2_decap_8 FILLER_62_1275 ();
 sg13g2_decap_8 FILLER_62_1282 ();
 sg13g2_decap_8 FILLER_62_1289 ();
 sg13g2_decap_8 FILLER_62_1296 ();
 sg13g2_decap_8 FILLER_62_1303 ();
 sg13g2_decap_4 FILLER_62_1310 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_11 ();
 sg13g2_decap_4 FILLER_63_18 ();
 sg13g2_fill_1 FILLER_63_22 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_106 ();
 sg13g2_fill_2 FILLER_63_143 ();
 sg13g2_fill_1 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_180 ();
 sg13g2_decap_4 FILLER_63_187 ();
 sg13g2_decap_8 FILLER_63_195 ();
 sg13g2_decap_8 FILLER_63_202 ();
 sg13g2_fill_2 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_215 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_4 FILLER_63_349 ();
 sg13g2_fill_1 FILLER_63_353 ();
 sg13g2_decap_8 FILLER_63_358 ();
 sg13g2_decap_4 FILLER_63_365 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_fill_1 FILLER_63_401 ();
 sg13g2_fill_2 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_63_410 ();
 sg13g2_decap_4 FILLER_63_431 ();
 sg13g2_fill_1 FILLER_63_435 ();
 sg13g2_fill_2 FILLER_63_442 ();
 sg13g2_fill_1 FILLER_63_444 ();
 sg13g2_decap_4 FILLER_63_449 ();
 sg13g2_fill_1 FILLER_63_453 ();
 sg13g2_fill_1 FILLER_63_482 ();
 sg13g2_fill_2 FILLER_63_496 ();
 sg13g2_decap_8 FILLER_63_506 ();
 sg13g2_fill_2 FILLER_63_513 ();
 sg13g2_decap_8 FILLER_63_561 ();
 sg13g2_decap_4 FILLER_63_568 ();
 sg13g2_fill_1 FILLER_63_572 ();
 sg13g2_fill_1 FILLER_63_621 ();
 sg13g2_decap_8 FILLER_63_647 ();
 sg13g2_decap_4 FILLER_63_654 ();
 sg13g2_decap_8 FILLER_63_662 ();
 sg13g2_fill_2 FILLER_63_669 ();
 sg13g2_fill_1 FILLER_63_671 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_fill_2 FILLER_63_714 ();
 sg13g2_fill_1 FILLER_63_716 ();
 sg13g2_decap_4 FILLER_63_740 ();
 sg13g2_decap_8 FILLER_63_748 ();
 sg13g2_fill_1 FILLER_63_755 ();
 sg13g2_decap_8 FILLER_63_760 ();
 sg13g2_decap_4 FILLER_63_767 ();
 sg13g2_fill_1 FILLER_63_771 ();
 sg13g2_decap_4 FILLER_63_785 ();
 sg13g2_fill_1 FILLER_63_793 ();
 sg13g2_decap_4 FILLER_63_804 ();
 sg13g2_fill_1 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_fill_1 FILLER_63_837 ();
 sg13g2_fill_2 FILLER_63_842 ();
 sg13g2_fill_1 FILLER_63_844 ();
 sg13g2_fill_2 FILLER_63_855 ();
 sg13g2_decap_8 FILLER_63_865 ();
 sg13g2_fill_2 FILLER_63_872 ();
 sg13g2_fill_1 FILLER_63_874 ();
 sg13g2_fill_1 FILLER_63_879 ();
 sg13g2_fill_2 FILLER_63_939 ();
 sg13g2_fill_1 FILLER_63_941 ();
 sg13g2_fill_1 FILLER_63_1046 ();
 sg13g2_fill_2 FILLER_63_1066 ();
 sg13g2_decap_8 FILLER_63_1104 ();
 sg13g2_decap_8 FILLER_63_1111 ();
 sg13g2_decap_8 FILLER_63_1118 ();
 sg13g2_decap_8 FILLER_63_1125 ();
 sg13g2_decap_8 FILLER_63_1132 ();
 sg13g2_decap_8 FILLER_63_1139 ();
 sg13g2_decap_8 FILLER_63_1146 ();
 sg13g2_decap_8 FILLER_63_1153 ();
 sg13g2_decap_8 FILLER_63_1160 ();
 sg13g2_decap_8 FILLER_63_1167 ();
 sg13g2_decap_8 FILLER_63_1174 ();
 sg13g2_decap_8 FILLER_63_1181 ();
 sg13g2_decap_8 FILLER_63_1188 ();
 sg13g2_decap_8 FILLER_63_1195 ();
 sg13g2_decap_8 FILLER_63_1202 ();
 sg13g2_decap_8 FILLER_63_1209 ();
 sg13g2_decap_8 FILLER_63_1216 ();
 sg13g2_decap_8 FILLER_63_1223 ();
 sg13g2_decap_8 FILLER_63_1230 ();
 sg13g2_decap_8 FILLER_63_1237 ();
 sg13g2_decap_8 FILLER_63_1244 ();
 sg13g2_decap_8 FILLER_63_1251 ();
 sg13g2_decap_8 FILLER_63_1258 ();
 sg13g2_decap_8 FILLER_63_1265 ();
 sg13g2_decap_8 FILLER_63_1272 ();
 sg13g2_decap_8 FILLER_63_1279 ();
 sg13g2_decap_8 FILLER_63_1286 ();
 sg13g2_decap_8 FILLER_63_1293 ();
 sg13g2_decap_8 FILLER_63_1300 ();
 sg13g2_decap_8 FILLER_63_1307 ();
 sg13g2_fill_1 FILLER_63_1314 ();
 sg13g2_decap_8 FILLER_64_26 ();
 sg13g2_decap_8 FILLER_64_33 ();
 sg13g2_decap_8 FILLER_64_40 ();
 sg13g2_fill_2 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_decap_4 FILLER_64_81 ();
 sg13g2_fill_2 FILLER_64_85 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_93 ();
 sg13g2_decap_8 FILLER_64_99 ();
 sg13g2_fill_1 FILLER_64_106 ();
 sg13g2_decap_4 FILLER_64_112 ();
 sg13g2_fill_1 FILLER_64_116 ();
 sg13g2_decap_4 FILLER_64_136 ();
 sg13g2_fill_1 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_145 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_fill_2 FILLER_64_159 ();
 sg13g2_fill_1 FILLER_64_161 ();
 sg13g2_decap_4 FILLER_64_214 ();
 sg13g2_decap_8 FILLER_64_222 ();
 sg13g2_fill_1 FILLER_64_229 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_2 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_269 ();
 sg13g2_fill_2 FILLER_64_280 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_fill_1 FILLER_64_366 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_decap_8 FILLER_64_436 ();
 sg13g2_decap_8 FILLER_64_443 ();
 sg13g2_decap_4 FILLER_64_450 ();
 sg13g2_fill_2 FILLER_64_454 ();
 sg13g2_decap_4 FILLER_64_468 ();
 sg13g2_fill_2 FILLER_64_477 ();
 sg13g2_fill_2 FILLER_64_491 ();
 sg13g2_fill_1 FILLER_64_493 ();
 sg13g2_decap_4 FILLER_64_512 ();
 sg13g2_fill_1 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_530 ();
 sg13g2_decap_8 FILLER_64_537 ();
 sg13g2_decap_8 FILLER_64_587 ();
 sg13g2_fill_2 FILLER_64_594 ();
 sg13g2_decap_8 FILLER_64_604 ();
 sg13g2_decap_4 FILLER_64_624 ();
 sg13g2_fill_1 FILLER_64_628 ();
 sg13g2_fill_2 FILLER_64_673 ();
 sg13g2_fill_1 FILLER_64_675 ();
 sg13g2_fill_2 FILLER_64_681 ();
 sg13g2_decap_8 FILLER_64_688 ();
 sg13g2_fill_2 FILLER_64_695 ();
 sg13g2_fill_1 FILLER_64_697 ();
 sg13g2_decap_4 FILLER_64_729 ();
 sg13g2_fill_2 FILLER_64_733 ();
 sg13g2_decap_4 FILLER_64_779 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_fill_2 FILLER_64_834 ();
 sg13g2_fill_1 FILLER_64_836 ();
 sg13g2_fill_2 FILLER_64_852 ();
 sg13g2_fill_2 FILLER_64_898 ();
 sg13g2_decap_8 FILLER_64_904 ();
 sg13g2_fill_1 FILLER_64_911 ();
 sg13g2_fill_2 FILLER_64_943 ();
 sg13g2_decap_8 FILLER_64_955 ();
 sg13g2_fill_2 FILLER_64_962 ();
 sg13g2_fill_2 FILLER_64_990 ();
 sg13g2_decap_8 FILLER_64_1009 ();
 sg13g2_fill_2 FILLER_64_1016 ();
 sg13g2_decap_4 FILLER_64_1022 ();
 sg13g2_fill_2 FILLER_64_1026 ();
 sg13g2_decap_4 FILLER_64_1037 ();
 sg13g2_fill_1 FILLER_64_1041 ();
 sg13g2_fill_2 FILLER_64_1065 ();
 sg13g2_decap_8 FILLER_64_1107 ();
 sg13g2_decap_8 FILLER_64_1114 ();
 sg13g2_decap_8 FILLER_64_1121 ();
 sg13g2_decap_8 FILLER_64_1128 ();
 sg13g2_decap_8 FILLER_64_1135 ();
 sg13g2_decap_8 FILLER_64_1142 ();
 sg13g2_decap_8 FILLER_64_1149 ();
 sg13g2_decap_8 FILLER_64_1156 ();
 sg13g2_decap_8 FILLER_64_1163 ();
 sg13g2_decap_8 FILLER_64_1170 ();
 sg13g2_decap_8 FILLER_64_1177 ();
 sg13g2_decap_8 FILLER_64_1184 ();
 sg13g2_decap_8 FILLER_64_1191 ();
 sg13g2_decap_8 FILLER_64_1198 ();
 sg13g2_decap_8 FILLER_64_1205 ();
 sg13g2_decap_8 FILLER_64_1212 ();
 sg13g2_decap_8 FILLER_64_1219 ();
 sg13g2_decap_8 FILLER_64_1226 ();
 sg13g2_decap_8 FILLER_64_1233 ();
 sg13g2_decap_8 FILLER_64_1240 ();
 sg13g2_decap_8 FILLER_64_1247 ();
 sg13g2_decap_8 FILLER_64_1254 ();
 sg13g2_decap_8 FILLER_64_1261 ();
 sg13g2_decap_8 FILLER_64_1268 ();
 sg13g2_decap_8 FILLER_64_1275 ();
 sg13g2_decap_8 FILLER_64_1282 ();
 sg13g2_decap_8 FILLER_64_1289 ();
 sg13g2_decap_8 FILLER_64_1296 ();
 sg13g2_decap_8 FILLER_64_1303 ();
 sg13g2_decap_4 FILLER_64_1310 ();
 sg13g2_fill_1 FILLER_64_1314 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_41 ();
 sg13g2_decap_4 FILLER_65_45 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_64 ();
 sg13g2_decap_8 FILLER_65_117 ();
 sg13g2_fill_1 FILLER_65_124 ();
 sg13g2_fill_2 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_132 ();
 sg13g2_decap_4 FILLER_65_171 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_2 FILLER_65_182 ();
 sg13g2_decap_4 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_192 ();
 sg13g2_fill_1 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_2 FILLER_65_313 ();
 sg13g2_fill_1 FILLER_65_315 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_338 ();
 sg13g2_decap_8 FILLER_65_345 ();
 sg13g2_decap_8 FILLER_65_352 ();
 sg13g2_fill_2 FILLER_65_359 ();
 sg13g2_decap_8 FILLER_65_365 ();
 sg13g2_decap_4 FILLER_65_372 ();
 sg13g2_fill_1 FILLER_65_376 ();
 sg13g2_fill_2 FILLER_65_388 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_4 FILLER_65_412 ();
 sg13g2_fill_2 FILLER_65_424 ();
 sg13g2_fill_1 FILLER_65_426 ();
 sg13g2_decap_4 FILLER_65_453 ();
 sg13g2_fill_1 FILLER_65_457 ();
 sg13g2_fill_1 FILLER_65_484 ();
 sg13g2_decap_4 FILLER_65_501 ();
 sg13g2_fill_2 FILLER_65_510 ();
 sg13g2_fill_1 FILLER_65_512 ();
 sg13g2_decap_4 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_553 ();
 sg13g2_decap_4 FILLER_65_559 ();
 sg13g2_fill_2 FILLER_65_563 ();
 sg13g2_fill_2 FILLER_65_626 ();
 sg13g2_fill_1 FILLER_65_628 ();
 sg13g2_fill_2 FILLER_65_633 ();
 sg13g2_decap_4 FILLER_65_645 ();
 sg13g2_fill_2 FILLER_65_649 ();
 sg13g2_decap_8 FILLER_65_659 ();
 sg13g2_decap_8 FILLER_65_666 ();
 sg13g2_fill_2 FILLER_65_673 ();
 sg13g2_fill_1 FILLER_65_675 ();
 sg13g2_decap_4 FILLER_65_681 ();
 sg13g2_fill_1 FILLER_65_708 ();
 sg13g2_decap_4 FILLER_65_761 ();
 sg13g2_decap_4 FILLER_65_773 ();
 sg13g2_fill_2 FILLER_65_777 ();
 sg13g2_fill_1 FILLER_65_792 ();
 sg13g2_decap_4 FILLER_65_807 ();
 sg13g2_fill_2 FILLER_65_811 ();
 sg13g2_fill_1 FILLER_65_843 ();
 sg13g2_fill_2 FILLER_65_895 ();
 sg13g2_decap_8 FILLER_65_923 ();
 sg13g2_fill_1 FILLER_65_930 ();
 sg13g2_decap_4 FILLER_65_957 ();
 sg13g2_decap_4 FILLER_65_971 ();
 sg13g2_decap_8 FILLER_65_979 ();
 sg13g2_decap_4 FILLER_65_986 ();
 sg13g2_decap_8 FILLER_65_993 ();
 sg13g2_decap_4 FILLER_65_1000 ();
 sg13g2_fill_1 FILLER_65_1004 ();
 sg13g2_decap_8 FILLER_65_1018 ();
 sg13g2_decap_8 FILLER_65_1057 ();
 sg13g2_fill_1 FILLER_65_1064 ();
 sg13g2_decap_8 FILLER_65_1075 ();
 sg13g2_fill_2 FILLER_65_1082 ();
 sg13g2_decap_8 FILLER_65_1101 ();
 sg13g2_decap_8 FILLER_65_1108 ();
 sg13g2_decap_8 FILLER_65_1115 ();
 sg13g2_decap_8 FILLER_65_1122 ();
 sg13g2_decap_8 FILLER_65_1129 ();
 sg13g2_decap_8 FILLER_65_1136 ();
 sg13g2_decap_8 FILLER_65_1143 ();
 sg13g2_decap_8 FILLER_65_1150 ();
 sg13g2_decap_8 FILLER_65_1157 ();
 sg13g2_decap_8 FILLER_65_1164 ();
 sg13g2_decap_8 FILLER_65_1171 ();
 sg13g2_decap_8 FILLER_65_1178 ();
 sg13g2_decap_8 FILLER_65_1185 ();
 sg13g2_decap_8 FILLER_65_1192 ();
 sg13g2_decap_8 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1206 ();
 sg13g2_decap_8 FILLER_65_1213 ();
 sg13g2_decap_8 FILLER_65_1220 ();
 sg13g2_decap_8 FILLER_65_1227 ();
 sg13g2_decap_8 FILLER_65_1234 ();
 sg13g2_decap_8 FILLER_65_1241 ();
 sg13g2_decap_8 FILLER_65_1248 ();
 sg13g2_decap_8 FILLER_65_1255 ();
 sg13g2_decap_8 FILLER_65_1262 ();
 sg13g2_decap_8 FILLER_65_1269 ();
 sg13g2_decap_8 FILLER_65_1276 ();
 sg13g2_decap_8 FILLER_65_1283 ();
 sg13g2_decap_8 FILLER_65_1290 ();
 sg13g2_decap_8 FILLER_65_1297 ();
 sg13g2_decap_8 FILLER_65_1304 ();
 sg13g2_decap_4 FILLER_65_1311 ();
 sg13g2_decap_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_2 FILLER_66_13 ();
 sg13g2_decap_4 FILLER_66_23 ();
 sg13g2_fill_2 FILLER_66_30 ();
 sg13g2_decap_4 FILLER_66_37 ();
 sg13g2_decap_8 FILLER_66_67 ();
 sg13g2_fill_2 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_76 ();
 sg13g2_fill_2 FILLER_66_85 ();
 sg13g2_fill_1 FILLER_66_87 ();
 sg13g2_fill_1 FILLER_66_94 ();
 sg13g2_fill_2 FILLER_66_109 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_fill_2 FILLER_66_164 ();
 sg13g2_decap_8 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_decap_8 FILLER_66_209 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_2 FILLER_66_326 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_decap_4 FILLER_66_338 ();
 sg13g2_fill_2 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_405 ();
 sg13g2_fill_2 FILLER_66_412 ();
 sg13g2_decap_8 FILLER_66_455 ();
 sg13g2_decap_8 FILLER_66_462 ();
 sg13g2_decap_8 FILLER_66_473 ();
 sg13g2_decap_4 FILLER_66_480 ();
 sg13g2_fill_1 FILLER_66_484 ();
 sg13g2_fill_2 FILLER_66_511 ();
 sg13g2_fill_1 FILLER_66_513 ();
 sg13g2_decap_4 FILLER_66_528 ();
 sg13g2_fill_2 FILLER_66_532 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_fill_1 FILLER_66_587 ();
 sg13g2_fill_2 FILLER_66_596 ();
 sg13g2_fill_1 FILLER_66_598 ();
 sg13g2_decap_8 FILLER_66_603 ();
 sg13g2_decap_4 FILLER_66_610 ();
 sg13g2_fill_1 FILLER_66_617 ();
 sg13g2_fill_2 FILLER_66_644 ();
 sg13g2_decap_8 FILLER_66_715 ();
 sg13g2_decap_4 FILLER_66_722 ();
 sg13g2_fill_2 FILLER_66_726 ();
 sg13g2_fill_2 FILLER_66_732 ();
 sg13g2_decap_4 FILLER_66_770 ();
 sg13g2_decap_8 FILLER_66_813 ();
 sg13g2_fill_2 FILLER_66_829 ();
 sg13g2_fill_1 FILLER_66_831 ();
 sg13g2_fill_2 FILLER_66_842 ();
 sg13g2_fill_1 FILLER_66_844 ();
 sg13g2_decap_4 FILLER_66_849 ();
 sg13g2_fill_2 FILLER_66_857 ();
 sg13g2_fill_1 FILLER_66_859 ();
 sg13g2_decap_8 FILLER_66_870 ();
 sg13g2_fill_2 FILLER_66_877 ();
 sg13g2_fill_1 FILLER_66_879 ();
 sg13g2_decap_4 FILLER_66_884 ();
 sg13g2_fill_1 FILLER_66_888 ();
 sg13g2_decap_8 FILLER_66_914 ();
 sg13g2_decap_8 FILLER_66_921 ();
 sg13g2_fill_2 FILLER_66_936 ();
 sg13g2_decap_8 FILLER_66_947 ();
 sg13g2_fill_1 FILLER_66_954 ();
 sg13g2_decap_8 FILLER_66_996 ();
 sg13g2_decap_4 FILLER_66_1043 ();
 sg13g2_fill_1 FILLER_66_1047 ();
 sg13g2_decap_8 FILLER_66_1100 ();
 sg13g2_decap_8 FILLER_66_1107 ();
 sg13g2_decap_8 FILLER_66_1114 ();
 sg13g2_decap_8 FILLER_66_1121 ();
 sg13g2_decap_8 FILLER_66_1128 ();
 sg13g2_decap_8 FILLER_66_1135 ();
 sg13g2_decap_8 FILLER_66_1142 ();
 sg13g2_decap_8 FILLER_66_1149 ();
 sg13g2_decap_8 FILLER_66_1156 ();
 sg13g2_decap_8 FILLER_66_1163 ();
 sg13g2_decap_8 FILLER_66_1170 ();
 sg13g2_decap_8 FILLER_66_1177 ();
 sg13g2_decap_8 FILLER_66_1184 ();
 sg13g2_decap_8 FILLER_66_1191 ();
 sg13g2_decap_8 FILLER_66_1198 ();
 sg13g2_decap_8 FILLER_66_1205 ();
 sg13g2_decap_8 FILLER_66_1212 ();
 sg13g2_decap_8 FILLER_66_1219 ();
 sg13g2_decap_8 FILLER_66_1226 ();
 sg13g2_decap_8 FILLER_66_1233 ();
 sg13g2_decap_8 FILLER_66_1240 ();
 sg13g2_decap_8 FILLER_66_1247 ();
 sg13g2_decap_8 FILLER_66_1254 ();
 sg13g2_decap_8 FILLER_66_1261 ();
 sg13g2_decap_8 FILLER_66_1268 ();
 sg13g2_decap_8 FILLER_66_1275 ();
 sg13g2_decap_8 FILLER_66_1282 ();
 sg13g2_decap_8 FILLER_66_1289 ();
 sg13g2_decap_8 FILLER_66_1296 ();
 sg13g2_decap_8 FILLER_66_1303 ();
 sg13g2_decap_4 FILLER_66_1310 ();
 sg13g2_fill_1 FILLER_66_1314 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_28 ();
 sg13g2_fill_1 FILLER_67_46 ();
 sg13g2_decap_8 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_101 ();
 sg13g2_decap_4 FILLER_67_110 ();
 sg13g2_decap_4 FILLER_67_117 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_133 ();
 sg13g2_fill_1 FILLER_67_135 ();
 sg13g2_decap_8 FILLER_67_150 ();
 sg13g2_fill_2 FILLER_67_157 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_2 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_185 ();
 sg13g2_fill_2 FILLER_67_192 ();
 sg13g2_decap_4 FILLER_67_200 ();
 sg13g2_fill_1 FILLER_67_204 ();
 sg13g2_fill_1 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_253 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_fill_2 FILLER_67_268 ();
 sg13g2_fill_1 FILLER_67_270 ();
 sg13g2_fill_2 FILLER_67_320 ();
 sg13g2_decap_8 FILLER_67_353 ();
 sg13g2_decap_4 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_377 ();
 sg13g2_fill_2 FILLER_67_419 ();
 sg13g2_fill_1 FILLER_67_421 ();
 sg13g2_decap_4 FILLER_67_433 ();
 sg13g2_fill_1 FILLER_67_437 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_fill_2 FILLER_67_545 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_fill_2 FILLER_67_552 ();
 sg13g2_fill_1 FILLER_67_554 ();
 sg13g2_fill_2 FILLER_67_559 ();
 sg13g2_fill_2 FILLER_67_565 ();
 sg13g2_fill_2 FILLER_67_585 ();
 sg13g2_fill_1 FILLER_67_587 ();
 sg13g2_decap_4 FILLER_67_629 ();
 sg13g2_decap_4 FILLER_67_638 ();
 sg13g2_fill_1 FILLER_67_642 ();
 sg13g2_fill_1 FILLER_67_658 ();
 sg13g2_decap_4 FILLER_67_669 ();
 sg13g2_fill_2 FILLER_67_677 ();
 sg13g2_fill_1 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_690 ();
 sg13g2_fill_2 FILLER_67_697 ();
 sg13g2_fill_1 FILLER_67_699 ();
 sg13g2_fill_1 FILLER_67_709 ();
 sg13g2_fill_2 FILLER_67_749 ();
 sg13g2_fill_1 FILLER_67_751 ();
 sg13g2_decap_8 FILLER_67_764 ();
 sg13g2_decap_8 FILLER_67_771 ();
 sg13g2_fill_1 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_789 ();
 sg13g2_fill_2 FILLER_67_796 ();
 sg13g2_fill_1 FILLER_67_798 ();
 sg13g2_fill_2 FILLER_67_811 ();
 sg13g2_fill_1 FILLER_67_813 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_fill_1 FILLER_67_878 ();
 sg13g2_decap_4 FILLER_67_883 ();
 sg13g2_fill_2 FILLER_67_887 ();
 sg13g2_decap_4 FILLER_67_910 ();
 sg13g2_fill_2 FILLER_67_914 ();
 sg13g2_decap_4 FILLER_67_968 ();
 sg13g2_decap_4 FILLER_67_977 ();
 sg13g2_fill_1 FILLER_67_985 ();
 sg13g2_fill_1 FILLER_67_993 ();
 sg13g2_decap_8 FILLER_67_1007 ();
 sg13g2_decap_4 FILLER_67_1018 ();
 sg13g2_fill_1 FILLER_67_1027 ();
 sg13g2_fill_1 FILLER_67_1033 ();
 sg13g2_decap_4 FILLER_67_1038 ();
 sg13g2_fill_2 FILLER_67_1050 ();
 sg13g2_decap_4 FILLER_67_1057 ();
 sg13g2_fill_1 FILLER_67_1061 ();
 sg13g2_decap_8 FILLER_67_1071 ();
 sg13g2_decap_8 FILLER_67_1078 ();
 sg13g2_decap_8 FILLER_67_1092 ();
 sg13g2_decap_8 FILLER_67_1099 ();
 sg13g2_decap_8 FILLER_67_1106 ();
 sg13g2_decap_8 FILLER_67_1113 ();
 sg13g2_decap_8 FILLER_67_1120 ();
 sg13g2_decap_8 FILLER_67_1127 ();
 sg13g2_decap_8 FILLER_67_1134 ();
 sg13g2_decap_8 FILLER_67_1141 ();
 sg13g2_decap_8 FILLER_67_1148 ();
 sg13g2_decap_8 FILLER_67_1155 ();
 sg13g2_decap_8 FILLER_67_1162 ();
 sg13g2_decap_8 FILLER_67_1169 ();
 sg13g2_decap_8 FILLER_67_1176 ();
 sg13g2_decap_8 FILLER_67_1183 ();
 sg13g2_decap_8 FILLER_67_1190 ();
 sg13g2_decap_8 FILLER_67_1197 ();
 sg13g2_decap_8 FILLER_67_1204 ();
 sg13g2_decap_8 FILLER_67_1211 ();
 sg13g2_decap_8 FILLER_67_1218 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_decap_8 FILLER_67_1232 ();
 sg13g2_decap_8 FILLER_67_1239 ();
 sg13g2_decap_8 FILLER_67_1246 ();
 sg13g2_decap_8 FILLER_67_1253 ();
 sg13g2_decap_8 FILLER_67_1260 ();
 sg13g2_decap_8 FILLER_67_1267 ();
 sg13g2_decap_8 FILLER_67_1274 ();
 sg13g2_decap_8 FILLER_67_1281 ();
 sg13g2_decap_8 FILLER_67_1288 ();
 sg13g2_decap_8 FILLER_67_1295 ();
 sg13g2_decap_8 FILLER_67_1302 ();
 sg13g2_decap_4 FILLER_67_1309 ();
 sg13g2_fill_2 FILLER_67_1313 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_35 ();
 sg13g2_fill_2 FILLER_68_50 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_decap_4 FILLER_68_65 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_222 ();
 sg13g2_fill_1 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_284 ();
 sg13g2_decap_4 FILLER_68_320 ();
 sg13g2_fill_1 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_decap_4 FILLER_68_377 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_398 ();
 sg13g2_fill_1 FILLER_68_451 ();
 sg13g2_decap_8 FILLER_68_499 ();
 sg13g2_fill_2 FILLER_68_506 ();
 sg13g2_decap_8 FILLER_68_512 ();
 sg13g2_decap_4 FILLER_68_519 ();
 sg13g2_fill_2 FILLER_68_523 ();
 sg13g2_decap_4 FILLER_68_546 ();
 sg13g2_fill_1 FILLER_68_550 ();
 sg13g2_decap_4 FILLER_68_587 ();
 sg13g2_fill_1 FILLER_68_591 ();
 sg13g2_decap_4 FILLER_68_602 ();
 sg13g2_fill_1 FILLER_68_606 ();
 sg13g2_fill_2 FILLER_68_617 ();
 sg13g2_fill_1 FILLER_68_619 ();
 sg13g2_fill_2 FILLER_68_636 ();
 sg13g2_decap_4 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_718 ();
 sg13g2_fill_1 FILLER_68_720 ();
 sg13g2_decap_4 FILLER_68_725 ();
 sg13g2_fill_1 FILLER_68_729 ();
 sg13g2_fill_1 FILLER_68_743 ();
 sg13g2_fill_1 FILLER_68_752 ();
 sg13g2_fill_1 FILLER_68_772 ();
 sg13g2_fill_1 FILLER_68_802 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_fill_2 FILLER_68_825 ();
 sg13g2_fill_1 FILLER_68_827 ();
 sg13g2_decap_8 FILLER_68_842 ();
 sg13g2_fill_1 FILLER_68_857 ();
 sg13g2_decap_8 FILLER_68_894 ();
 sg13g2_decap_8 FILLER_68_901 ();
 sg13g2_fill_1 FILLER_68_908 ();
 sg13g2_fill_2 FILLER_68_917 ();
 sg13g2_fill_1 FILLER_68_919 ();
 sg13g2_decap_8 FILLER_68_939 ();
 sg13g2_fill_2 FILLER_68_946 ();
 sg13g2_fill_1 FILLER_68_948 ();
 sg13g2_decap_4 FILLER_68_958 ();
 sg13g2_fill_2 FILLER_68_962 ();
 sg13g2_fill_2 FILLER_68_983 ();
 sg13g2_fill_2 FILLER_68_1008 ();
 sg13g2_fill_1 FILLER_68_1010 ();
 sg13g2_fill_2 FILLER_68_1016 ();
 sg13g2_fill_1 FILLER_68_1018 ();
 sg13g2_fill_2 FILLER_68_1027 ();
 sg13g2_fill_1 FILLER_68_1029 ();
 sg13g2_fill_1 FILLER_68_1049 ();
 sg13g2_decap_4 FILLER_68_1063 ();
 sg13g2_fill_1 FILLER_68_1067 ();
 sg13g2_decap_8 FILLER_68_1104 ();
 sg13g2_decap_8 FILLER_68_1111 ();
 sg13g2_decap_8 FILLER_68_1118 ();
 sg13g2_decap_8 FILLER_68_1125 ();
 sg13g2_decap_8 FILLER_68_1132 ();
 sg13g2_decap_8 FILLER_68_1139 ();
 sg13g2_decap_8 FILLER_68_1146 ();
 sg13g2_decap_8 FILLER_68_1153 ();
 sg13g2_decap_8 FILLER_68_1160 ();
 sg13g2_decap_8 FILLER_68_1167 ();
 sg13g2_decap_8 FILLER_68_1174 ();
 sg13g2_decap_8 FILLER_68_1181 ();
 sg13g2_decap_8 FILLER_68_1188 ();
 sg13g2_decap_8 FILLER_68_1195 ();
 sg13g2_decap_8 FILLER_68_1202 ();
 sg13g2_decap_8 FILLER_68_1209 ();
 sg13g2_decap_8 FILLER_68_1216 ();
 sg13g2_decap_8 FILLER_68_1223 ();
 sg13g2_decap_8 FILLER_68_1230 ();
 sg13g2_decap_8 FILLER_68_1237 ();
 sg13g2_decap_8 FILLER_68_1244 ();
 sg13g2_decap_8 FILLER_68_1251 ();
 sg13g2_decap_8 FILLER_68_1258 ();
 sg13g2_decap_8 FILLER_68_1265 ();
 sg13g2_decap_8 FILLER_68_1272 ();
 sg13g2_decap_8 FILLER_68_1279 ();
 sg13g2_decap_8 FILLER_68_1286 ();
 sg13g2_decap_8 FILLER_68_1293 ();
 sg13g2_decap_8 FILLER_68_1300 ();
 sg13g2_decap_8 FILLER_68_1307 ();
 sg13g2_fill_1 FILLER_68_1314 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_17 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_4 FILLER_69_169 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_decap_8 FILLER_69_179 ();
 sg13g2_fill_2 FILLER_69_189 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_2 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_242 ();
 sg13g2_decap_4 FILLER_69_249 ();
 sg13g2_fill_2 FILLER_69_253 ();
 sg13g2_decap_4 FILLER_69_262 ();
 sg13g2_fill_2 FILLER_69_266 ();
 sg13g2_fill_2 FILLER_69_280 ();
 sg13g2_fill_2 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_288 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_4 FILLER_69_308 ();
 sg13g2_fill_1 FILLER_69_345 ();
 sg13g2_decap_8 FILLER_69_354 ();
 sg13g2_fill_1 FILLER_69_361 ();
 sg13g2_decap_4 FILLER_69_366 ();
 sg13g2_fill_2 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_fill_2 FILLER_69_397 ();
 sg13g2_decap_8 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_410 ();
 sg13g2_decap_8 FILLER_69_422 ();
 sg13g2_decap_4 FILLER_69_429 ();
 sg13g2_fill_1 FILLER_69_433 ();
 sg13g2_fill_2 FILLER_69_442 ();
 sg13g2_decap_8 FILLER_69_454 ();
 sg13g2_fill_2 FILLER_69_461 ();
 sg13g2_fill_1 FILLER_69_467 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_fill_2 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_538 ();
 sg13g2_decap_8 FILLER_69_545 ();
 sg13g2_fill_2 FILLER_69_552 ();
 sg13g2_fill_1 FILLER_69_554 ();
 sg13g2_decap_8 FILLER_69_559 ();
 sg13g2_decap_4 FILLER_69_566 ();
 sg13g2_fill_1 FILLER_69_570 ();
 sg13g2_fill_2 FILLER_69_580 ();
 sg13g2_fill_1 FILLER_69_586 ();
 sg13g2_fill_1 FILLER_69_630 ();
 sg13g2_decap_4 FILLER_69_636 ();
 sg13g2_fill_1 FILLER_69_640 ();
 sg13g2_decap_8 FILLER_69_648 ();
 sg13g2_decap_4 FILLER_69_655 ();
 sg13g2_fill_2 FILLER_69_669 ();
 sg13g2_fill_1 FILLER_69_671 ();
 sg13g2_fill_2 FILLER_69_676 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_decap_8 FILLER_69_689 ();
 sg13g2_decap_4 FILLER_69_696 ();
 sg13g2_fill_2 FILLER_69_726 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_742 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_fill_1 FILLER_69_756 ();
 sg13g2_decap_4 FILLER_69_762 ();
 sg13g2_fill_2 FILLER_69_781 ();
 sg13g2_fill_1 FILLER_69_783 ();
 sg13g2_decap_8 FILLER_69_788 ();
 sg13g2_decap_4 FILLER_69_795 ();
 sg13g2_fill_2 FILLER_69_799 ();
 sg13g2_fill_2 FILLER_69_819 ();
 sg13g2_decap_4 FILLER_69_847 ();
 sg13g2_fill_1 FILLER_69_851 ();
 sg13g2_decap_8 FILLER_69_885 ();
 sg13g2_fill_1 FILLER_69_892 ();
 sg13g2_fill_2 FILLER_69_943 ();
 sg13g2_fill_1 FILLER_69_945 ();
 sg13g2_decap_4 FILLER_69_959 ();
 sg13g2_fill_1 FILLER_69_963 ();
 sg13g2_decap_4 FILLER_69_967 ();
 sg13g2_fill_2 FILLER_69_991 ();
 sg13g2_decap_4 FILLER_69_1005 ();
 sg13g2_decap_4 FILLER_69_1017 ();
 sg13g2_fill_1 FILLER_69_1021 ();
 sg13g2_decap_8 FILLER_69_1026 ();
 sg13g2_fill_2 FILLER_69_1049 ();
 sg13g2_fill_1 FILLER_69_1051 ();
 sg13g2_decap_8 FILLER_69_1065 ();
 sg13g2_decap_8 FILLER_69_1072 ();
 sg13g2_decap_8 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1094 ();
 sg13g2_decap_8 FILLER_69_1101 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_decap_8 FILLER_69_1115 ();
 sg13g2_decap_8 FILLER_69_1122 ();
 sg13g2_decap_8 FILLER_69_1129 ();
 sg13g2_decap_8 FILLER_69_1136 ();
 sg13g2_decap_8 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1157 ();
 sg13g2_decap_8 FILLER_69_1164 ();
 sg13g2_decap_8 FILLER_69_1171 ();
 sg13g2_decap_8 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1185 ();
 sg13g2_decap_8 FILLER_69_1192 ();
 sg13g2_decap_8 FILLER_69_1199 ();
 sg13g2_decap_8 FILLER_69_1206 ();
 sg13g2_decap_8 FILLER_69_1213 ();
 sg13g2_decap_8 FILLER_69_1220 ();
 sg13g2_decap_8 FILLER_69_1227 ();
 sg13g2_decap_8 FILLER_69_1234 ();
 sg13g2_decap_8 FILLER_69_1241 ();
 sg13g2_decap_8 FILLER_69_1248 ();
 sg13g2_decap_8 FILLER_69_1255 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_decap_8 FILLER_69_1269 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_decap_8 FILLER_69_1283 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_4 FILLER_69_1311 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_33 ();
 sg13g2_decap_8 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_44 ();
 sg13g2_fill_1 FILLER_70_46 ();
 sg13g2_decap_8 FILLER_70_50 ();
 sg13g2_decap_8 FILLER_70_57 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_82 ();
 sg13g2_fill_1 FILLER_70_84 ();
 sg13g2_decap_4 FILLER_70_90 ();
 sg13g2_fill_2 FILLER_70_94 ();
 sg13g2_fill_2 FILLER_70_114 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_1 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_2 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_236 ();
 sg13g2_decap_4 FILLER_70_248 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_258 ();
 sg13g2_fill_1 FILLER_70_265 ();
 sg13g2_fill_2 FILLER_70_271 ();
 sg13g2_decap_4 FILLER_70_289 ();
 sg13g2_decap_4 FILLER_70_310 ();
 sg13g2_fill_2 FILLER_70_314 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_322 ();
 sg13g2_fill_1 FILLER_70_327 ();
 sg13g2_decap_8 FILLER_70_375 ();
 sg13g2_decap_8 FILLER_70_382 ();
 sg13g2_decap_4 FILLER_70_415 ();
 sg13g2_fill_2 FILLER_70_419 ();
 sg13g2_fill_2 FILLER_70_447 ();
 sg13g2_decap_4 FILLER_70_492 ();
 sg13g2_decap_8 FILLER_70_500 ();
 sg13g2_fill_2 FILLER_70_507 ();
 sg13g2_fill_1 FILLER_70_509 ();
 sg13g2_decap_8 FILLER_70_536 ();
 sg13g2_fill_1 FILLER_70_543 ();
 sg13g2_fill_2 FILLER_70_580 ();
 sg13g2_decap_8 FILLER_70_605 ();
 sg13g2_fill_2 FILLER_70_612 ();
 sg13g2_fill_1 FILLER_70_632 ();
 sg13g2_decap_4 FILLER_70_638 ();
 sg13g2_decap_8 FILLER_70_650 ();
 sg13g2_fill_2 FILLER_70_657 ();
 sg13g2_fill_2 FILLER_70_671 ();
 sg13g2_decap_8 FILLER_70_677 ();
 sg13g2_fill_2 FILLER_70_684 ();
 sg13g2_decap_4 FILLER_70_691 ();
 sg13g2_fill_1 FILLER_70_710 ();
 sg13g2_decap_8 FILLER_70_715 ();
 sg13g2_fill_1 FILLER_70_722 ();
 sg13g2_fill_2 FILLER_70_726 ();
 sg13g2_fill_1 FILLER_70_728 ();
 sg13g2_decap_4 FILLER_70_742 ();
 sg13g2_fill_2 FILLER_70_746 ();
 sg13g2_fill_2 FILLER_70_754 ();
 sg13g2_fill_1 FILLER_70_756 ();
 sg13g2_fill_1 FILLER_70_816 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_fill_2 FILLER_70_829 ();
 sg13g2_fill_1 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_836 ();
 sg13g2_decap_4 FILLER_70_843 ();
 sg13g2_fill_1 FILLER_70_853 ();
 sg13g2_decap_4 FILLER_70_899 ();
 sg13g2_fill_2 FILLER_70_928 ();
 sg13g2_fill_1 FILLER_70_966 ();
 sg13g2_fill_1 FILLER_70_989 ();
 sg13g2_fill_1 FILLER_70_1037 ();
 sg13g2_fill_2 FILLER_70_1041 ();
 sg13g2_decap_4 FILLER_70_1061 ();
 sg13g2_fill_1 FILLER_70_1065 ();
 sg13g2_decap_8 FILLER_70_1102 ();
 sg13g2_decap_8 FILLER_70_1109 ();
 sg13g2_decap_8 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_decap_8 FILLER_70_1137 ();
 sg13g2_decap_8 FILLER_70_1144 ();
 sg13g2_decap_8 FILLER_70_1151 ();
 sg13g2_decap_8 FILLER_70_1158 ();
 sg13g2_decap_8 FILLER_70_1165 ();
 sg13g2_decap_8 FILLER_70_1172 ();
 sg13g2_decap_8 FILLER_70_1179 ();
 sg13g2_decap_8 FILLER_70_1186 ();
 sg13g2_decap_8 FILLER_70_1193 ();
 sg13g2_decap_8 FILLER_70_1200 ();
 sg13g2_decap_8 FILLER_70_1207 ();
 sg13g2_decap_8 FILLER_70_1214 ();
 sg13g2_decap_8 FILLER_70_1221 ();
 sg13g2_decap_8 FILLER_70_1228 ();
 sg13g2_decap_8 FILLER_70_1235 ();
 sg13g2_decap_8 FILLER_70_1242 ();
 sg13g2_decap_8 FILLER_70_1249 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1263 ();
 sg13g2_decap_8 FILLER_70_1270 ();
 sg13g2_decap_8 FILLER_70_1277 ();
 sg13g2_decap_8 FILLER_70_1284 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_8 FILLER_70_1298 ();
 sg13g2_decap_8 FILLER_70_1305 ();
 sg13g2_fill_2 FILLER_70_1312 ();
 sg13g2_fill_1 FILLER_70_1314 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_4 ();
 sg13g2_fill_2 FILLER_71_9 ();
 sg13g2_fill_1 FILLER_71_11 ();
 sg13g2_fill_2 FILLER_71_48 ();
 sg13g2_fill_1 FILLER_71_50 ();
 sg13g2_decap_4 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_69 ();
 sg13g2_decap_8 FILLER_71_75 ();
 sg13g2_fill_2 FILLER_71_82 ();
 sg13g2_fill_1 FILLER_71_84 ();
 sg13g2_fill_2 FILLER_71_101 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_147 ();
 sg13g2_decap_4 FILLER_71_158 ();
 sg13g2_decap_8 FILLER_71_166 ();
 sg13g2_fill_2 FILLER_71_173 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_decap_4 FILLER_71_199 ();
 sg13g2_decap_8 FILLER_71_212 ();
 sg13g2_fill_2 FILLER_71_219 ();
 sg13g2_fill_2 FILLER_71_225 ();
 sg13g2_fill_2 FILLER_71_232 ();
 sg13g2_fill_1 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_368 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_2 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_fill_2 FILLER_71_421 ();
 sg13g2_fill_1 FILLER_71_423 ();
 sg13g2_fill_2 FILLER_71_428 ();
 sg13g2_fill_1 FILLER_71_430 ();
 sg13g2_decap_8 FILLER_71_435 ();
 sg13g2_fill_2 FILLER_71_442 ();
 sg13g2_decap_4 FILLER_71_454 ();
 sg13g2_fill_2 FILLER_71_458 ();
 sg13g2_decap_8 FILLER_71_464 ();
 sg13g2_fill_2 FILLER_71_471 ();
 sg13g2_fill_1 FILLER_71_473 ();
 sg13g2_decap_8 FILLER_71_500 ();
 sg13g2_decap_4 FILLER_71_507 ();
 sg13g2_fill_1 FILLER_71_511 ();
 sg13g2_fill_2 FILLER_71_526 ();
 sg13g2_decap_4 FILLER_71_564 ();
 sg13g2_fill_1 FILLER_71_568 ();
 sg13g2_decap_8 FILLER_71_588 ();
 sg13g2_decap_8 FILLER_71_595 ();
 sg13g2_fill_1 FILLER_71_602 ();
 sg13g2_decap_4 FILLER_71_628 ();
 sg13g2_fill_2 FILLER_71_650 ();
 sg13g2_fill_1 FILLER_71_720 ();
 sg13g2_fill_1 FILLER_71_725 ();
 sg13g2_fill_1 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_775 ();
 sg13g2_decap_4 FILLER_71_782 ();
 sg13g2_decap_4 FILLER_71_790 ();
 sg13g2_fill_2 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_fill_2 FILLER_71_831 ();
 sg13g2_fill_1 FILLER_71_833 ();
 sg13g2_fill_1 FILLER_71_860 ();
 sg13g2_decap_4 FILLER_71_869 ();
 sg13g2_decap_8 FILLER_71_913 ();
 sg13g2_fill_1 FILLER_71_920 ();
 sg13g2_decap_4 FILLER_71_934 ();
 sg13g2_fill_2 FILLER_71_948 ();
 sg13g2_fill_1 FILLER_71_950 ();
 sg13g2_decap_8 FILLER_71_955 ();
 sg13g2_decap_4 FILLER_71_962 ();
 sg13g2_fill_1 FILLER_71_966 ();
 sg13g2_fill_1 FILLER_71_977 ();
 sg13g2_fill_1 FILLER_71_988 ();
 sg13g2_decap_8 FILLER_71_994 ();
 sg13g2_fill_1 FILLER_71_1001 ();
 sg13g2_decap_4 FILLER_71_1012 ();
 sg13g2_fill_2 FILLER_71_1016 ();
 sg13g2_decap_8 FILLER_71_1022 ();
 sg13g2_decap_8 FILLER_71_1029 ();
 sg13g2_fill_2 FILLER_71_1036 ();
 sg13g2_fill_1 FILLER_71_1051 ();
 sg13g2_fill_2 FILLER_71_1055 ();
 sg13g2_decap_8 FILLER_71_1083 ();
 sg13g2_decap_8 FILLER_71_1090 ();
 sg13g2_decap_8 FILLER_71_1097 ();
 sg13g2_decap_8 FILLER_71_1104 ();
 sg13g2_decap_8 FILLER_71_1111 ();
 sg13g2_decap_8 FILLER_71_1118 ();
 sg13g2_decap_8 FILLER_71_1125 ();
 sg13g2_decap_8 FILLER_71_1132 ();
 sg13g2_decap_8 FILLER_71_1139 ();
 sg13g2_decap_8 FILLER_71_1146 ();
 sg13g2_decap_8 FILLER_71_1153 ();
 sg13g2_decap_8 FILLER_71_1160 ();
 sg13g2_decap_8 FILLER_71_1167 ();
 sg13g2_decap_8 FILLER_71_1174 ();
 sg13g2_decap_8 FILLER_71_1181 ();
 sg13g2_decap_8 FILLER_71_1188 ();
 sg13g2_decap_8 FILLER_71_1195 ();
 sg13g2_decap_8 FILLER_71_1202 ();
 sg13g2_decap_8 FILLER_71_1209 ();
 sg13g2_decap_8 FILLER_71_1216 ();
 sg13g2_decap_8 FILLER_71_1223 ();
 sg13g2_decap_8 FILLER_71_1230 ();
 sg13g2_decap_8 FILLER_71_1237 ();
 sg13g2_decap_8 FILLER_71_1244 ();
 sg13g2_decap_8 FILLER_71_1251 ();
 sg13g2_decap_8 FILLER_71_1258 ();
 sg13g2_decap_8 FILLER_71_1265 ();
 sg13g2_decap_8 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1293 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_fill_1 FILLER_71_1314 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_17 ();
 sg13g2_decap_4 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_34 ();
 sg13g2_decap_4 FILLER_72_39 ();
 sg13g2_fill_2 FILLER_72_127 ();
 sg13g2_fill_1 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_140 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_decap_4 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_1 FILLER_72_249 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_decap_4 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_290 ();
 sg13g2_fill_2 FILLER_72_302 ();
 sg13g2_fill_1 FILLER_72_304 ();
 sg13g2_fill_1 FILLER_72_310 ();
 sg13g2_fill_1 FILLER_72_320 ();
 sg13g2_fill_2 FILLER_72_347 ();
 sg13g2_decap_8 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_360 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_2 FILLER_72_379 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_fill_1 FILLER_72_387 ();
 sg13g2_decap_4 FILLER_72_440 ();
 sg13g2_fill_1 FILLER_72_444 ();
 sg13g2_fill_1 FILLER_72_497 ();
 sg13g2_fill_2 FILLER_72_545 ();
 sg13g2_fill_1 FILLER_72_547 ();
 sg13g2_fill_2 FILLER_72_552 ();
 sg13g2_fill_2 FILLER_72_587 ();
 sg13g2_fill_1 FILLER_72_589 ();
 sg13g2_fill_2 FILLER_72_616 ();
 sg13g2_fill_1 FILLER_72_618 ();
 sg13g2_fill_2 FILLER_72_627 ();
 sg13g2_decap_4 FILLER_72_635 ();
 sg13g2_decap_4 FILLER_72_649 ();
 sg13g2_decap_4 FILLER_72_661 ();
 sg13g2_fill_2 FILLER_72_692 ();
 sg13g2_fill_1 FILLER_72_694 ();
 sg13g2_decap_4 FILLER_72_742 ();
 sg13g2_fill_2 FILLER_72_784 ();
 sg13g2_fill_1 FILLER_72_786 ();
 sg13g2_decap_4 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_800 ();
 sg13g2_decap_4 FILLER_72_854 ();
 sg13g2_fill_1 FILLER_72_858 ();
 sg13g2_fill_1 FILLER_72_863 ();
 sg13g2_fill_2 FILLER_72_872 ();
 sg13g2_fill_1 FILLER_72_874 ();
 sg13g2_decap_8 FILLER_72_901 ();
 sg13g2_decap_8 FILLER_72_908 ();
 sg13g2_decap_4 FILLER_72_915 ();
 sg13g2_fill_1 FILLER_72_945 ();
 sg13g2_decap_4 FILLER_72_977 ();
 sg13g2_fill_2 FILLER_72_1007 ();
 sg13g2_fill_1 FILLER_72_1009 ();
 sg13g2_fill_2 FILLER_72_1062 ();
 sg13g2_fill_1 FILLER_72_1064 ();
 sg13g2_decap_8 FILLER_72_1079 ();
 sg13g2_decap_8 FILLER_72_1086 ();
 sg13g2_decap_8 FILLER_72_1093 ();
 sg13g2_decap_8 FILLER_72_1100 ();
 sg13g2_decap_8 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_decap_8 FILLER_72_1121 ();
 sg13g2_decap_8 FILLER_72_1128 ();
 sg13g2_decap_8 FILLER_72_1135 ();
 sg13g2_decap_8 FILLER_72_1142 ();
 sg13g2_decap_8 FILLER_72_1149 ();
 sg13g2_decap_8 FILLER_72_1156 ();
 sg13g2_decap_8 FILLER_72_1163 ();
 sg13g2_decap_8 FILLER_72_1170 ();
 sg13g2_decap_8 FILLER_72_1177 ();
 sg13g2_decap_8 FILLER_72_1184 ();
 sg13g2_decap_8 FILLER_72_1191 ();
 sg13g2_decap_8 FILLER_72_1198 ();
 sg13g2_decap_8 FILLER_72_1205 ();
 sg13g2_decap_8 FILLER_72_1212 ();
 sg13g2_decap_8 FILLER_72_1219 ();
 sg13g2_decap_8 FILLER_72_1226 ();
 sg13g2_decap_8 FILLER_72_1233 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_decap_8 FILLER_72_1247 ();
 sg13g2_decap_8 FILLER_72_1254 ();
 sg13g2_decap_8 FILLER_72_1261 ();
 sg13g2_decap_8 FILLER_72_1268 ();
 sg13g2_decap_8 FILLER_72_1275 ();
 sg13g2_decap_8 FILLER_72_1282 ();
 sg13g2_decap_8 FILLER_72_1289 ();
 sg13g2_decap_8 FILLER_72_1296 ();
 sg13g2_decap_8 FILLER_72_1303 ();
 sg13g2_decap_4 FILLER_72_1310 ();
 sg13g2_fill_1 FILLER_72_1314 ();
 sg13g2_fill_1 FILLER_73_26 ();
 sg13g2_fill_2 FILLER_73_35 ();
 sg13g2_fill_1 FILLER_73_37 ();
 sg13g2_fill_1 FILLER_73_48 ();
 sg13g2_decap_4 FILLER_73_65 ();
 sg13g2_decap_8 FILLER_73_72 ();
 sg13g2_decap_8 FILLER_73_83 ();
 sg13g2_decap_4 FILLER_73_90 ();
 sg13g2_fill_1 FILLER_73_94 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_fill_2 FILLER_73_105 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_decap_4 FILLER_73_172 ();
 sg13g2_fill_1 FILLER_73_176 ();
 sg13g2_fill_2 FILLER_73_191 ();
 sg13g2_decap_8 FILLER_73_198 ();
 sg13g2_decap_4 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_decap_8 FILLER_73_290 ();
 sg13g2_fill_2 FILLER_73_307 ();
 sg13g2_decap_4 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_378 ();
 sg13g2_fill_1 FILLER_73_380 ();
 sg13g2_decap_4 FILLER_73_385 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_fill_2 FILLER_73_401 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_73_414 ();
 sg13g2_fill_2 FILLER_73_457 ();
 sg13g2_fill_1 FILLER_73_459 ();
 sg13g2_decap_4 FILLER_73_464 ();
 sg13g2_decap_4 FILLER_73_478 ();
 sg13g2_fill_2 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_488 ();
 sg13g2_decap_4 FILLER_73_519 ();
 sg13g2_fill_1 FILLER_73_523 ();
 sg13g2_decap_8 FILLER_73_545 ();
 sg13g2_decap_8 FILLER_73_552 ();
 sg13g2_decap_8 FILLER_73_559 ();
 sg13g2_decap_4 FILLER_73_566 ();
 sg13g2_fill_1 FILLER_73_570 ();
 sg13g2_decap_8 FILLER_73_586 ();
 sg13g2_decap_4 FILLER_73_593 ();
 sg13g2_decap_8 FILLER_73_611 ();
 sg13g2_fill_1 FILLER_73_626 ();
 sg13g2_decap_4 FILLER_73_658 ();
 sg13g2_fill_2 FILLER_73_662 ();
 sg13g2_fill_2 FILLER_73_685 ();
 sg13g2_fill_1 FILLER_73_687 ();
 sg13g2_fill_2 FILLER_73_701 ();
 sg13g2_fill_1 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_decap_4 FILLER_73_716 ();
 sg13g2_fill_1 FILLER_73_720 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_fill_1 FILLER_73_814 ();
 sg13g2_fill_2 FILLER_73_866 ();
 sg13g2_decap_8 FILLER_73_878 ();
 sg13g2_fill_1 FILLER_73_885 ();
 sg13g2_decap_4 FILLER_73_916 ();
 sg13g2_fill_1 FILLER_73_920 ();
 sg13g2_decap_8 FILLER_73_947 ();
 sg13g2_fill_1 FILLER_73_954 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_fill_1 FILLER_73_976 ();
 sg13g2_decap_4 FILLER_73_987 ();
 sg13g2_fill_1 FILLER_73_991 ();
 sg13g2_decap_4 FILLER_73_996 ();
 sg13g2_decap_8 FILLER_73_1003 ();
 sg13g2_decap_4 FILLER_73_1010 ();
 sg13g2_fill_1 FILLER_73_1014 ();
 sg13g2_fill_1 FILLER_73_1029 ();
 sg13g2_decap_8 FILLER_73_1034 ();
 sg13g2_decap_4 FILLER_73_1041 ();
 sg13g2_fill_1 FILLER_73_1045 ();
 sg13g2_fill_2 FILLER_73_1050 ();
 sg13g2_fill_1 FILLER_73_1052 ();
 sg13g2_decap_8 FILLER_73_1063 ();
 sg13g2_decap_8 FILLER_73_1070 ();
 sg13g2_decap_8 FILLER_73_1077 ();
 sg13g2_decap_8 FILLER_73_1084 ();
 sg13g2_decap_8 FILLER_73_1091 ();
 sg13g2_decap_8 FILLER_73_1098 ();
 sg13g2_decap_8 FILLER_73_1105 ();
 sg13g2_decap_8 FILLER_73_1112 ();
 sg13g2_decap_8 FILLER_73_1119 ();
 sg13g2_decap_8 FILLER_73_1126 ();
 sg13g2_decap_8 FILLER_73_1133 ();
 sg13g2_decap_8 FILLER_73_1140 ();
 sg13g2_decap_8 FILLER_73_1147 ();
 sg13g2_decap_8 FILLER_73_1154 ();
 sg13g2_decap_8 FILLER_73_1161 ();
 sg13g2_decap_8 FILLER_73_1168 ();
 sg13g2_decap_8 FILLER_73_1175 ();
 sg13g2_decap_8 FILLER_73_1182 ();
 sg13g2_decap_8 FILLER_73_1189 ();
 sg13g2_decap_8 FILLER_73_1196 ();
 sg13g2_decap_8 FILLER_73_1203 ();
 sg13g2_decap_8 FILLER_73_1210 ();
 sg13g2_decap_8 FILLER_73_1217 ();
 sg13g2_decap_8 FILLER_73_1224 ();
 sg13g2_decap_8 FILLER_73_1231 ();
 sg13g2_decap_8 FILLER_73_1238 ();
 sg13g2_decap_8 FILLER_73_1245 ();
 sg13g2_decap_8 FILLER_73_1252 ();
 sg13g2_decap_8 FILLER_73_1259 ();
 sg13g2_decap_8 FILLER_73_1266 ();
 sg13g2_decap_8 FILLER_73_1273 ();
 sg13g2_decap_8 FILLER_73_1280 ();
 sg13g2_decap_8 FILLER_73_1287 ();
 sg13g2_decap_8 FILLER_73_1294 ();
 sg13g2_decap_8 FILLER_73_1301 ();
 sg13g2_decap_8 FILLER_73_1308 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_15 ();
 sg13g2_fill_1 FILLER_74_25 ();
 sg13g2_fill_2 FILLER_74_30 ();
 sg13g2_fill_2 FILLER_74_47 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_fill_2 FILLER_74_128 ();
 sg13g2_fill_2 FILLER_74_143 ();
 sg13g2_decap_8 FILLER_74_149 ();
 sg13g2_fill_2 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_158 ();
 sg13g2_fill_2 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_250 ();
 sg13g2_decap_4 FILLER_74_255 ();
 sg13g2_fill_2 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_307 ();
 sg13g2_fill_2 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_316 ();
 sg13g2_decap_4 FILLER_74_342 ();
 sg13g2_fill_1 FILLER_74_346 ();
 sg13g2_fill_2 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_421 ();
 sg13g2_decap_4 FILLER_74_428 ();
 sg13g2_fill_1 FILLER_74_432 ();
 sg13g2_decap_4 FILLER_74_441 ();
 sg13g2_decap_4 FILLER_74_454 ();
 sg13g2_decap_8 FILLER_74_466 ();
 sg13g2_decap_8 FILLER_74_473 ();
 sg13g2_decap_8 FILLER_74_480 ();
 sg13g2_decap_8 FILLER_74_487 ();
 sg13g2_decap_4 FILLER_74_494 ();
 sg13g2_fill_2 FILLER_74_498 ();
 sg13g2_fill_1 FILLER_74_504 ();
 sg13g2_decap_8 FILLER_74_520 ();
 sg13g2_fill_2 FILLER_74_527 ();
 sg13g2_fill_1 FILLER_74_529 ();
 sg13g2_decap_4 FILLER_74_540 ();
 sg13g2_decap_4 FILLER_74_569 ();
 sg13g2_fill_1 FILLER_74_573 ();
 sg13g2_fill_2 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_628 ();
 sg13g2_fill_2 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_640 ();
 sg13g2_fill_2 FILLER_74_647 ();
 sg13g2_fill_1 FILLER_74_649 ();
 sg13g2_fill_2 FILLER_74_686 ();
 sg13g2_fill_1 FILLER_74_688 ();
 sg13g2_fill_2 FILLER_74_699 ();
 sg13g2_fill_2 FILLER_74_758 ();
 sg13g2_decap_4 FILLER_74_764 ();
 sg13g2_fill_2 FILLER_74_768 ();
 sg13g2_decap_4 FILLER_74_790 ();
 sg13g2_fill_1 FILLER_74_794 ();
 sg13g2_fill_2 FILLER_74_799 ();
 sg13g2_fill_2 FILLER_74_811 ();
 sg13g2_decap_4 FILLER_74_826 ();
 sg13g2_fill_1 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_845 ();
 sg13g2_decap_4 FILLER_74_870 ();
 sg13g2_fill_2 FILLER_74_874 ();
 sg13g2_fill_2 FILLER_74_902 ();
 sg13g2_fill_1 FILLER_74_904 ();
 sg13g2_fill_1 FILLER_74_931 ();
 sg13g2_fill_2 FILLER_74_941 ();
 sg13g2_fill_1 FILLER_74_943 ();
 sg13g2_decap_4 FILLER_74_952 ();
 sg13g2_fill_1 FILLER_74_982 ();
 sg13g2_decap_8 FILLER_74_1009 ();
 sg13g2_fill_2 FILLER_74_1016 ();
 sg13g2_fill_1 FILLER_74_1018 ();
 sg13g2_decap_8 FILLER_74_1045 ();
 sg13g2_decap_8 FILLER_74_1052 ();
 sg13g2_decap_8 FILLER_74_1059 ();
 sg13g2_decap_8 FILLER_74_1066 ();
 sg13g2_decap_8 FILLER_74_1073 ();
 sg13g2_decap_8 FILLER_74_1080 ();
 sg13g2_decap_8 FILLER_74_1087 ();
 sg13g2_decap_8 FILLER_74_1094 ();
 sg13g2_decap_8 FILLER_74_1101 ();
 sg13g2_decap_8 FILLER_74_1108 ();
 sg13g2_decap_8 FILLER_74_1115 ();
 sg13g2_decap_8 FILLER_74_1122 ();
 sg13g2_decap_8 FILLER_74_1129 ();
 sg13g2_decap_8 FILLER_74_1136 ();
 sg13g2_decap_8 FILLER_74_1143 ();
 sg13g2_decap_8 FILLER_74_1150 ();
 sg13g2_decap_8 FILLER_74_1157 ();
 sg13g2_decap_8 FILLER_74_1164 ();
 sg13g2_decap_8 FILLER_74_1171 ();
 sg13g2_decap_8 FILLER_74_1178 ();
 sg13g2_decap_8 FILLER_74_1185 ();
 sg13g2_decap_8 FILLER_74_1192 ();
 sg13g2_decap_8 FILLER_74_1199 ();
 sg13g2_decap_8 FILLER_74_1206 ();
 sg13g2_decap_8 FILLER_74_1213 ();
 sg13g2_decap_8 FILLER_74_1220 ();
 sg13g2_decap_8 FILLER_74_1227 ();
 sg13g2_decap_8 FILLER_74_1234 ();
 sg13g2_decap_8 FILLER_74_1241 ();
 sg13g2_decap_8 FILLER_74_1248 ();
 sg13g2_decap_8 FILLER_74_1255 ();
 sg13g2_decap_8 FILLER_74_1262 ();
 sg13g2_decap_8 FILLER_74_1269 ();
 sg13g2_decap_8 FILLER_74_1276 ();
 sg13g2_decap_8 FILLER_74_1283 ();
 sg13g2_decap_8 FILLER_74_1290 ();
 sg13g2_decap_8 FILLER_74_1297 ();
 sg13g2_decap_8 FILLER_74_1304 ();
 sg13g2_decap_4 FILLER_74_1311 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_16 ();
 sg13g2_fill_1 FILLER_75_47 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_2 FILLER_75_145 ();
 sg13g2_fill_2 FILLER_75_151 ();
 sg13g2_fill_2 FILLER_75_173 ();
 sg13g2_fill_2 FILLER_75_178 ();
 sg13g2_decap_8 FILLER_75_188 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_197 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_4 FILLER_75_231 ();
 sg13g2_fill_2 FILLER_75_235 ();
 sg13g2_fill_2 FILLER_75_247 ();
 sg13g2_decap_4 FILLER_75_269 ();
 sg13g2_fill_2 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_353 ();
 sg13g2_fill_2 FILLER_75_370 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_fill_2 FILLER_75_428 ();
 sg13g2_fill_1 FILLER_75_456 ();
 sg13g2_fill_1 FILLER_75_466 ();
 sg13g2_decap_4 FILLER_75_503 ();
 sg13g2_fill_1 FILLER_75_507 ();
 sg13g2_fill_2 FILLER_75_581 ();
 sg13g2_fill_1 FILLER_75_583 ();
 sg13g2_fill_2 FILLER_75_588 ();
 sg13g2_fill_1 FILLER_75_590 ();
 sg13g2_decap_8 FILLER_75_601 ();
 sg13g2_decap_4 FILLER_75_634 ();
 sg13g2_decap_8 FILLER_75_648 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_fill_2 FILLER_75_671 ();
 sg13g2_fill_1 FILLER_75_673 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_fill_2 FILLER_75_712 ();
 sg13g2_fill_1 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_4 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_4 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_870 ();
 sg13g2_decap_8 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_75_884 ();
 sg13g2_fill_1 FILLER_75_886 ();
 sg13g2_decap_8 FILLER_75_891 ();
 sg13g2_decap_4 FILLER_75_898 ();
 sg13g2_fill_2 FILLER_75_912 ();
 sg13g2_fill_1 FILLER_75_914 ();
 sg13g2_decap_8 FILLER_75_919 ();
 sg13g2_decap_4 FILLER_75_926 ();
 sg13g2_fill_1 FILLER_75_930 ();
 sg13g2_decap_4 FILLER_75_935 ();
 sg13g2_fill_1 FILLER_75_939 ();
 sg13g2_fill_2 FILLER_75_950 ();
 sg13g2_decap_8 FILLER_75_957 ();
 sg13g2_fill_2 FILLER_75_964 ();
 sg13g2_fill_1 FILLER_75_966 ();
 sg13g2_decap_8 FILLER_75_971 ();
 sg13g2_decap_8 FILLER_75_978 ();
 sg13g2_decap_8 FILLER_75_985 ();
 sg13g2_fill_2 FILLER_75_992 ();
 sg13g2_decap_8 FILLER_75_998 ();
 sg13g2_decap_8 FILLER_75_1005 ();
 sg13g2_decap_8 FILLER_75_1012 ();
 sg13g2_decap_8 FILLER_75_1019 ();
 sg13g2_decap_8 FILLER_75_1026 ();
 sg13g2_decap_8 FILLER_75_1033 ();
 sg13g2_decap_8 FILLER_75_1040 ();
 sg13g2_decap_8 FILLER_75_1047 ();
 sg13g2_decap_8 FILLER_75_1054 ();
 sg13g2_decap_8 FILLER_75_1061 ();
 sg13g2_decap_8 FILLER_75_1068 ();
 sg13g2_decap_8 FILLER_75_1075 ();
 sg13g2_decap_8 FILLER_75_1082 ();
 sg13g2_decap_8 FILLER_75_1089 ();
 sg13g2_decap_8 FILLER_75_1096 ();
 sg13g2_decap_8 FILLER_75_1103 ();
 sg13g2_decap_8 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1117 ();
 sg13g2_decap_8 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1131 ();
 sg13g2_decap_8 FILLER_75_1138 ();
 sg13g2_decap_8 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1152 ();
 sg13g2_decap_8 FILLER_75_1159 ();
 sg13g2_decap_8 FILLER_75_1166 ();
 sg13g2_decap_8 FILLER_75_1173 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_decap_8 FILLER_75_1187 ();
 sg13g2_decap_8 FILLER_75_1194 ();
 sg13g2_decap_8 FILLER_75_1201 ();
 sg13g2_decap_8 FILLER_75_1208 ();
 sg13g2_decap_8 FILLER_75_1215 ();
 sg13g2_decap_8 FILLER_75_1222 ();
 sg13g2_decap_8 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1236 ();
 sg13g2_decap_8 FILLER_75_1243 ();
 sg13g2_decap_8 FILLER_75_1250 ();
 sg13g2_decap_8 FILLER_75_1257 ();
 sg13g2_decap_8 FILLER_75_1264 ();
 sg13g2_decap_8 FILLER_75_1271 ();
 sg13g2_decap_8 FILLER_75_1278 ();
 sg13g2_decap_8 FILLER_75_1285 ();
 sg13g2_decap_8 FILLER_75_1292 ();
 sg13g2_decap_8 FILLER_75_1299 ();
 sg13g2_decap_8 FILLER_75_1306 ();
 sg13g2_fill_2 FILLER_75_1313 ();
 sg13g2_fill_1 FILLER_76_26 ();
 sg13g2_fill_1 FILLER_76_37 ();
 sg13g2_fill_2 FILLER_76_47 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_4 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_81 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_decap_4 FILLER_76_109 ();
 sg13g2_fill_1 FILLER_76_113 ();
 sg13g2_fill_2 FILLER_76_145 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_235 ();
 sg13g2_fill_2 FILLER_76_250 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_fill_2 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_fill_1 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_324 ();
 sg13g2_fill_2 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_4 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_396 ();
 sg13g2_fill_1 FILLER_76_407 ();
 sg13g2_decap_4 FILLER_76_469 ();
 sg13g2_fill_2 FILLER_76_519 ();
 sg13g2_fill_1 FILLER_76_521 ();
 sg13g2_decap_8 FILLER_76_526 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_fill_2 FILLER_76_540 ();
 sg13g2_fill_1 FILLER_76_542 ();
 sg13g2_fill_2 FILLER_76_569 ();
 sg13g2_fill_2 FILLER_76_575 ();
 sg13g2_decap_8 FILLER_76_587 ();
 sg13g2_decap_4 FILLER_76_594 ();
 sg13g2_decap_4 FILLER_76_608 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_fill_2 FILLER_76_617 ();
 sg13g2_fill_2 FILLER_76_623 ();
 sg13g2_fill_2 FILLER_76_687 ();
 sg13g2_decap_4 FILLER_76_756 ();
 sg13g2_fill_2 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_fill_1 FILLER_76_777 ();
 sg13g2_decap_4 FILLER_76_793 ();
 sg13g2_fill_2 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_803 ();
 sg13g2_decap_8 FILLER_76_810 ();
 sg13g2_decap_8 FILLER_76_817 ();
 sg13g2_decap_4 FILLER_76_824 ();
 sg13g2_fill_2 FILLER_76_832 ();
 sg13g2_fill_1 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_845 ();
 sg13g2_fill_2 FILLER_76_852 ();
 sg13g2_fill_1 FILLER_76_854 ();
 sg13g2_fill_2 FILLER_76_859 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_fill_1 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_883 ();
 sg13g2_fill_2 FILLER_76_921 ();
 sg13g2_fill_1 FILLER_76_923 ();
 sg13g2_decap_8 FILLER_76_928 ();
 sg13g2_decap_8 FILLER_76_935 ();
 sg13g2_decap_8 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_949 ();
 sg13g2_decap_8 FILLER_76_956 ();
 sg13g2_decap_8 FILLER_76_963 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_decap_8 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_984 ();
 sg13g2_decap_8 FILLER_76_991 ();
 sg13g2_decap_8 FILLER_76_998 ();
 sg13g2_decap_8 FILLER_76_1005 ();
 sg13g2_decap_8 FILLER_76_1012 ();
 sg13g2_decap_8 FILLER_76_1019 ();
 sg13g2_decap_8 FILLER_76_1026 ();
 sg13g2_decap_8 FILLER_76_1033 ();
 sg13g2_decap_8 FILLER_76_1040 ();
 sg13g2_decap_8 FILLER_76_1047 ();
 sg13g2_decap_8 FILLER_76_1054 ();
 sg13g2_decap_8 FILLER_76_1061 ();
 sg13g2_decap_8 FILLER_76_1068 ();
 sg13g2_decap_8 FILLER_76_1075 ();
 sg13g2_decap_8 FILLER_76_1082 ();
 sg13g2_decap_8 FILLER_76_1089 ();
 sg13g2_decap_8 FILLER_76_1096 ();
 sg13g2_decap_8 FILLER_76_1103 ();
 sg13g2_decap_8 FILLER_76_1110 ();
 sg13g2_decap_8 FILLER_76_1117 ();
 sg13g2_decap_8 FILLER_76_1124 ();
 sg13g2_decap_8 FILLER_76_1131 ();
 sg13g2_decap_8 FILLER_76_1138 ();
 sg13g2_decap_8 FILLER_76_1145 ();
 sg13g2_decap_8 FILLER_76_1152 ();
 sg13g2_decap_8 FILLER_76_1159 ();
 sg13g2_decap_8 FILLER_76_1166 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_decap_8 FILLER_76_1180 ();
 sg13g2_decap_8 FILLER_76_1187 ();
 sg13g2_decap_8 FILLER_76_1194 ();
 sg13g2_decap_8 FILLER_76_1201 ();
 sg13g2_decap_8 FILLER_76_1208 ();
 sg13g2_decap_8 FILLER_76_1215 ();
 sg13g2_decap_8 FILLER_76_1222 ();
 sg13g2_decap_8 FILLER_76_1229 ();
 sg13g2_decap_8 FILLER_76_1236 ();
 sg13g2_decap_8 FILLER_76_1243 ();
 sg13g2_decap_8 FILLER_76_1250 ();
 sg13g2_decap_8 FILLER_76_1257 ();
 sg13g2_decap_8 FILLER_76_1264 ();
 sg13g2_decap_8 FILLER_76_1271 ();
 sg13g2_decap_8 FILLER_76_1278 ();
 sg13g2_decap_8 FILLER_76_1285 ();
 sg13g2_decap_8 FILLER_76_1292 ();
 sg13g2_decap_8 FILLER_76_1299 ();
 sg13g2_decap_8 FILLER_76_1306 ();
 sg13g2_fill_2 FILLER_76_1313 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_4 ();
 sg13g2_fill_1 FILLER_77_53 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_decap_4 FILLER_77_123 ();
 sg13g2_fill_2 FILLER_77_127 ();
 sg13g2_decap_8 FILLER_77_139 ();
 sg13g2_decap_4 FILLER_77_146 ();
 sg13g2_decap_4 FILLER_77_159 ();
 sg13g2_decap_4 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_249 ();
 sg13g2_decap_4 FILLER_77_254 ();
 sg13g2_decap_8 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_297 ();
 sg13g2_fill_2 FILLER_77_303 ();
 sg13g2_fill_1 FILLER_77_305 ();
 sg13g2_decap_8 FILLER_77_316 ();
 sg13g2_decap_4 FILLER_77_326 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_decap_8 FILLER_77_335 ();
 sg13g2_decap_8 FILLER_77_345 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_decap_4 FILLER_77_358 ();
 sg13g2_fill_1 FILLER_77_362 ();
 sg13g2_fill_2 FILLER_77_368 ();
 sg13g2_fill_1 FILLER_77_370 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_2 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_406 ();
 sg13g2_fill_2 FILLER_77_413 ();
 sg13g2_fill_2 FILLER_77_430 ();
 sg13g2_fill_1 FILLER_77_432 ();
 sg13g2_decap_8 FILLER_77_437 ();
 sg13g2_decap_8 FILLER_77_444 ();
 sg13g2_decap_8 FILLER_77_451 ();
 sg13g2_fill_2 FILLER_77_458 ();
 sg13g2_fill_1 FILLER_77_460 ();
 sg13g2_fill_1 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_480 ();
 sg13g2_fill_1 FILLER_77_487 ();
 sg13g2_fill_2 FILLER_77_492 ();
 sg13g2_decap_8 FILLER_77_498 ();
 sg13g2_fill_1 FILLER_77_505 ();
 sg13g2_fill_2 FILLER_77_552 ();
 sg13g2_fill_2 FILLER_77_558 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_4 FILLER_77_623 ();
 sg13g2_fill_1 FILLER_77_627 ();
 sg13g2_fill_2 FILLER_77_638 ();
 sg13g2_decap_8 FILLER_77_644 ();
 sg13g2_decap_8 FILLER_77_651 ();
 sg13g2_decap_4 FILLER_77_658 ();
 sg13g2_fill_2 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_fill_1 FILLER_77_707 ();
 sg13g2_decap_4 FILLER_77_713 ();
 sg13g2_fill_1 FILLER_77_717 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_fill_2 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_fill_2 FILLER_77_748 ();
 sg13g2_fill_2 FILLER_77_786 ();
 sg13g2_fill_1 FILLER_77_788 ();
 sg13g2_decap_4 FILLER_77_815 ();
 sg13g2_decap_4 FILLER_77_871 ();
 sg13g2_fill_2 FILLER_77_875 ();
 sg13g2_fill_2 FILLER_77_911 ();
 sg13g2_decap_8 FILLER_77_949 ();
 sg13g2_decap_8 FILLER_77_956 ();
 sg13g2_decap_8 FILLER_77_963 ();
 sg13g2_decap_8 FILLER_77_970 ();
 sg13g2_decap_8 FILLER_77_977 ();
 sg13g2_decap_8 FILLER_77_984 ();
 sg13g2_decap_8 FILLER_77_991 ();
 sg13g2_decap_8 FILLER_77_998 ();
 sg13g2_decap_8 FILLER_77_1005 ();
 sg13g2_decap_8 FILLER_77_1012 ();
 sg13g2_decap_8 FILLER_77_1019 ();
 sg13g2_decap_8 FILLER_77_1026 ();
 sg13g2_decap_8 FILLER_77_1033 ();
 sg13g2_decap_8 FILLER_77_1040 ();
 sg13g2_decap_8 FILLER_77_1047 ();
 sg13g2_decap_8 FILLER_77_1054 ();
 sg13g2_decap_8 FILLER_77_1061 ();
 sg13g2_decap_8 FILLER_77_1068 ();
 sg13g2_decap_8 FILLER_77_1075 ();
 sg13g2_decap_8 FILLER_77_1082 ();
 sg13g2_decap_8 FILLER_77_1089 ();
 sg13g2_decap_8 FILLER_77_1096 ();
 sg13g2_decap_8 FILLER_77_1103 ();
 sg13g2_decap_8 FILLER_77_1110 ();
 sg13g2_decap_8 FILLER_77_1117 ();
 sg13g2_decap_8 FILLER_77_1124 ();
 sg13g2_decap_8 FILLER_77_1131 ();
 sg13g2_decap_8 FILLER_77_1138 ();
 sg13g2_decap_8 FILLER_77_1145 ();
 sg13g2_decap_8 FILLER_77_1152 ();
 sg13g2_decap_8 FILLER_77_1159 ();
 sg13g2_decap_8 FILLER_77_1166 ();
 sg13g2_decap_8 FILLER_77_1173 ();
 sg13g2_decap_8 FILLER_77_1180 ();
 sg13g2_decap_8 FILLER_77_1187 ();
 sg13g2_decap_8 FILLER_77_1194 ();
 sg13g2_decap_8 FILLER_77_1201 ();
 sg13g2_decap_8 FILLER_77_1208 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_8 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1292 ();
 sg13g2_decap_8 FILLER_77_1299 ();
 sg13g2_decap_8 FILLER_77_1306 ();
 sg13g2_fill_2 FILLER_77_1313 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_11 ();
 sg13g2_fill_1 FILLER_78_30 ();
 sg13g2_fill_2 FILLER_78_79 ();
 sg13g2_fill_1 FILLER_78_81 ();
 sg13g2_fill_2 FILLER_78_99 ();
 sg13g2_fill_2 FILLER_78_127 ();
 sg13g2_decap_4 FILLER_78_166 ();
 sg13g2_fill_2 FILLER_78_170 ();
 sg13g2_decap_4 FILLER_78_180 ();
 sg13g2_decap_4 FILLER_78_214 ();
 sg13g2_fill_1 FILLER_78_218 ();
 sg13g2_decap_4 FILLER_78_239 ();
 sg13g2_decap_4 FILLER_78_276 ();
 sg13g2_fill_1 FILLER_78_280 ();
 sg13g2_fill_2 FILLER_78_299 ();
 sg13g2_decap_4 FILLER_78_327 ();
 sg13g2_fill_1 FILLER_78_331 ();
 sg13g2_fill_2 FILLER_78_394 ();
 sg13g2_decap_4 FILLER_78_409 ();
 sg13g2_decap_4 FILLER_78_432 ();
 sg13g2_fill_1 FILLER_78_436 ();
 sg13g2_fill_2 FILLER_78_471 ();
 sg13g2_fill_1 FILLER_78_473 ();
 sg13g2_decap_4 FILLER_78_504 ();
 sg13g2_fill_1 FILLER_78_508 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_4 FILLER_78_566 ();
 sg13g2_fill_2 FILLER_78_570 ();
 sg13g2_decap_8 FILLER_78_582 ();
 sg13g2_decap_4 FILLER_78_589 ();
 sg13g2_decap_8 FILLER_78_608 ();
 sg13g2_decap_8 FILLER_78_641 ();
 sg13g2_fill_1 FILLER_78_648 ();
 sg13g2_fill_1 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_712 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_fill_2 FILLER_78_752 ();
 sg13g2_decap_4 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_823 ();
 sg13g2_fill_2 FILLER_78_834 ();
 sg13g2_fill_1 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_fill_2 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_78_881 ();
 sg13g2_decap_8 FILLER_78_940 ();
 sg13g2_decap_8 FILLER_78_947 ();
 sg13g2_decap_8 FILLER_78_954 ();
 sg13g2_decap_8 FILLER_78_961 ();
 sg13g2_decap_8 FILLER_78_968 ();
 sg13g2_decap_8 FILLER_78_975 ();
 sg13g2_decap_8 FILLER_78_982 ();
 sg13g2_decap_8 FILLER_78_989 ();
 sg13g2_decap_8 FILLER_78_996 ();
 sg13g2_decap_8 FILLER_78_1003 ();
 sg13g2_decap_8 FILLER_78_1010 ();
 sg13g2_decap_8 FILLER_78_1017 ();
 sg13g2_decap_8 FILLER_78_1024 ();
 sg13g2_decap_8 FILLER_78_1031 ();
 sg13g2_decap_8 FILLER_78_1038 ();
 sg13g2_decap_8 FILLER_78_1045 ();
 sg13g2_decap_8 FILLER_78_1052 ();
 sg13g2_decap_8 FILLER_78_1059 ();
 sg13g2_decap_8 FILLER_78_1066 ();
 sg13g2_decap_8 FILLER_78_1073 ();
 sg13g2_decap_8 FILLER_78_1080 ();
 sg13g2_decap_8 FILLER_78_1087 ();
 sg13g2_decap_8 FILLER_78_1094 ();
 sg13g2_decap_8 FILLER_78_1101 ();
 sg13g2_decap_8 FILLER_78_1108 ();
 sg13g2_decap_8 FILLER_78_1115 ();
 sg13g2_decap_8 FILLER_78_1122 ();
 sg13g2_decap_8 FILLER_78_1129 ();
 sg13g2_decap_8 FILLER_78_1136 ();
 sg13g2_decap_8 FILLER_78_1143 ();
 sg13g2_decap_8 FILLER_78_1150 ();
 sg13g2_decap_8 FILLER_78_1157 ();
 sg13g2_decap_8 FILLER_78_1164 ();
 sg13g2_decap_8 FILLER_78_1171 ();
 sg13g2_decap_8 FILLER_78_1178 ();
 sg13g2_decap_8 FILLER_78_1185 ();
 sg13g2_decap_8 FILLER_78_1192 ();
 sg13g2_decap_8 FILLER_78_1199 ();
 sg13g2_decap_8 FILLER_78_1206 ();
 sg13g2_decap_8 FILLER_78_1213 ();
 sg13g2_decap_8 FILLER_78_1220 ();
 sg13g2_decap_8 FILLER_78_1227 ();
 sg13g2_decap_8 FILLER_78_1234 ();
 sg13g2_decap_8 FILLER_78_1241 ();
 sg13g2_decap_8 FILLER_78_1248 ();
 sg13g2_decap_8 FILLER_78_1255 ();
 sg13g2_decap_8 FILLER_78_1262 ();
 sg13g2_decap_8 FILLER_78_1269 ();
 sg13g2_decap_8 FILLER_78_1276 ();
 sg13g2_decap_8 FILLER_78_1283 ();
 sg13g2_decap_8 FILLER_78_1290 ();
 sg13g2_decap_8 FILLER_78_1297 ();
 sg13g2_decap_8 FILLER_78_1304 ();
 sg13g2_decap_4 FILLER_78_1311 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_4 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_52 ();
 sg13g2_decap_4 FILLER_79_83 ();
 sg13g2_fill_2 FILLER_79_87 ();
 sg13g2_decap_4 FILLER_79_122 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_135 ();
 sg13g2_fill_1 FILLER_79_142 ();
 sg13g2_decap_4 FILLER_79_147 ();
 sg13g2_fill_2 FILLER_79_164 ();
 sg13g2_fill_1 FILLER_79_166 ();
 sg13g2_decap_8 FILLER_79_171 ();
 sg13g2_decap_4 FILLER_79_178 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_fill_2 FILLER_79_196 ();
 sg13g2_fill_1 FILLER_79_198 ();
 sg13g2_fill_2 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_266 ();
 sg13g2_fill_2 FILLER_79_310 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_fill_2 FILLER_79_373 ();
 sg13g2_fill_1 FILLER_79_375 ();
 sg13g2_decap_4 FILLER_79_381 ();
 sg13g2_fill_2 FILLER_79_385 ();
 sg13g2_fill_2 FILLER_79_404 ();
 sg13g2_fill_2 FILLER_79_418 ();
 sg13g2_decap_4 FILLER_79_461 ();
 sg13g2_fill_1 FILLER_79_465 ();
 sg13g2_decap_4 FILLER_79_476 ();
 sg13g2_fill_2 FILLER_79_480 ();
 sg13g2_fill_1 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_fill_1 FILLER_79_546 ();
 sg13g2_fill_1 FILLER_79_625 ();
 sg13g2_fill_2 FILLER_79_630 ();
 sg13g2_fill_1 FILLER_79_632 ();
 sg13g2_decap_8 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_4 FILLER_79_675 ();
 sg13g2_decap_4 FILLER_79_725 ();
 sg13g2_fill_1 FILLER_79_729 ();
 sg13g2_fill_2 FILLER_79_738 ();
 sg13g2_decap_4 FILLER_79_786 ();
 sg13g2_fill_1 FILLER_79_790 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_fill_1 FILLER_79_876 ();
 sg13g2_fill_2 FILLER_79_903 ();
 sg13g2_decap_4 FILLER_79_915 ();
 sg13g2_fill_2 FILLER_79_919 ();
 sg13g2_fill_2 FILLER_79_925 ();
 sg13g2_fill_1 FILLER_79_927 ();
 sg13g2_decap_8 FILLER_79_938 ();
 sg13g2_decap_8 FILLER_79_945 ();
 sg13g2_decap_8 FILLER_79_952 ();
 sg13g2_decap_8 FILLER_79_959 ();
 sg13g2_decap_8 FILLER_79_966 ();
 sg13g2_decap_8 FILLER_79_973 ();
 sg13g2_decap_8 FILLER_79_980 ();
 sg13g2_decap_8 FILLER_79_987 ();
 sg13g2_decap_8 FILLER_79_994 ();
 sg13g2_decap_8 FILLER_79_1001 ();
 sg13g2_decap_8 FILLER_79_1008 ();
 sg13g2_decap_8 FILLER_79_1015 ();
 sg13g2_decap_8 FILLER_79_1022 ();
 sg13g2_decap_8 FILLER_79_1029 ();
 sg13g2_decap_8 FILLER_79_1036 ();
 sg13g2_decap_8 FILLER_79_1043 ();
 sg13g2_decap_8 FILLER_79_1050 ();
 sg13g2_decap_8 FILLER_79_1057 ();
 sg13g2_decap_8 FILLER_79_1064 ();
 sg13g2_decap_8 FILLER_79_1071 ();
 sg13g2_decap_8 FILLER_79_1078 ();
 sg13g2_decap_8 FILLER_79_1085 ();
 sg13g2_decap_8 FILLER_79_1092 ();
 sg13g2_decap_8 FILLER_79_1099 ();
 sg13g2_decap_8 FILLER_79_1106 ();
 sg13g2_decap_8 FILLER_79_1113 ();
 sg13g2_decap_8 FILLER_79_1120 ();
 sg13g2_decap_8 FILLER_79_1127 ();
 sg13g2_decap_8 FILLER_79_1134 ();
 sg13g2_decap_8 FILLER_79_1141 ();
 sg13g2_decap_8 FILLER_79_1148 ();
 sg13g2_decap_8 FILLER_79_1155 ();
 sg13g2_decap_8 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1169 ();
 sg13g2_decap_8 FILLER_79_1176 ();
 sg13g2_decap_8 FILLER_79_1183 ();
 sg13g2_decap_8 FILLER_79_1190 ();
 sg13g2_decap_8 FILLER_79_1197 ();
 sg13g2_decap_8 FILLER_79_1204 ();
 sg13g2_decap_8 FILLER_79_1211 ();
 sg13g2_decap_8 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1225 ();
 sg13g2_decap_8 FILLER_79_1232 ();
 sg13g2_decap_8 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1246 ();
 sg13g2_decap_8 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1260 ();
 sg13g2_decap_8 FILLER_79_1267 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_4 FILLER_79_1309 ();
 sg13g2_fill_2 FILLER_79_1313 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_9 ();
 sg13g2_fill_2 FILLER_80_36 ();
 sg13g2_decap_8 FILLER_80_41 ();
 sg13g2_decap_8 FILLER_80_48 ();
 sg13g2_fill_2 FILLER_80_58 ();
 sg13g2_fill_1 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_69 ();
 sg13g2_decap_8 FILLER_80_76 ();
 sg13g2_decap_8 FILLER_80_83 ();
 sg13g2_decap_8 FILLER_80_90 ();
 sg13g2_decap_4 FILLER_80_97 ();
 sg13g2_fill_2 FILLER_80_101 ();
 sg13g2_decap_8 FILLER_80_107 ();
 sg13g2_decap_4 FILLER_80_114 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_decap_8 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_146 ();
 sg13g2_fill_2 FILLER_80_153 ();
 sg13g2_fill_1 FILLER_80_155 ();
 sg13g2_decap_8 FILLER_80_182 ();
 sg13g2_decap_4 FILLER_80_189 ();
 sg13g2_fill_2 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_decap_8 FILLER_80_224 ();
 sg13g2_decap_4 FILLER_80_234 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_260 ();
 sg13g2_fill_2 FILLER_80_333 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_408 ();
 sg13g2_decap_4 FILLER_80_415 ();
 sg13g2_decap_4 FILLER_80_431 ();
 sg13g2_fill_1 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_fill_2 FILLER_80_469 ();
 sg13g2_decap_4 FILLER_80_497 ();
 sg13g2_fill_1 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_506 ();
 sg13g2_decap_4 FILLER_80_513 ();
 sg13g2_fill_2 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_fill_2 FILLER_80_535 ();
 sg13g2_decap_4 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_555 ();
 sg13g2_fill_2 FILLER_80_562 ();
 sg13g2_fill_1 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_569 ();
 sg13g2_decap_8 FILLER_80_576 ();
 sg13g2_fill_1 FILLER_80_583 ();
 sg13g2_fill_1 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_4 FILLER_80_606 ();
 sg13g2_decap_4 FILLER_80_614 ();
 sg13g2_fill_2 FILLER_80_648 ();
 sg13g2_fill_1 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_687 ();
 sg13g2_decap_4 FILLER_80_694 ();
 sg13g2_fill_1 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_703 ();
 sg13g2_fill_2 FILLER_80_710 ();
 sg13g2_fill_1 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_4 FILLER_80_756 ();
 sg13g2_fill_1 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_fill_2 FILLER_80_783 ();
 sg13g2_decap_4 FILLER_80_795 ();
 sg13g2_fill_2 FILLER_80_799 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_4 FILLER_80_830 ();
 sg13g2_fill_1 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_fill_2 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_859 ();
 sg13g2_decap_8 FILLER_80_866 ();
 sg13g2_decap_8 FILLER_80_873 ();
 sg13g2_decap_8 FILLER_80_880 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_fill_1 FILLER_80_898 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1036 ();
 sg13g2_decap_8 FILLER_80_1043 ();
 sg13g2_decap_8 FILLER_80_1050 ();
 sg13g2_decap_8 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_decap_8 FILLER_80_1071 ();
 sg13g2_decap_8 FILLER_80_1078 ();
 sg13g2_decap_8 FILLER_80_1085 ();
 sg13g2_decap_8 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1106 ();
 sg13g2_decap_8 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_decap_8 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1134 ();
 sg13g2_decap_8 FILLER_80_1141 ();
 sg13g2_decap_8 FILLER_80_1148 ();
 sg13g2_decap_8 FILLER_80_1155 ();
 sg13g2_decap_8 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1169 ();
 sg13g2_decap_8 FILLER_80_1176 ();
 sg13g2_decap_8 FILLER_80_1183 ();
 sg13g2_decap_8 FILLER_80_1190 ();
 sg13g2_decap_8 FILLER_80_1197 ();
 sg13g2_decap_8 FILLER_80_1204 ();
 sg13g2_decap_8 FILLER_80_1211 ();
 sg13g2_decap_8 FILLER_80_1218 ();
 sg13g2_decap_8 FILLER_80_1225 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_8 FILLER_80_1239 ();
 sg13g2_decap_8 FILLER_80_1246 ();
 sg13g2_decap_8 FILLER_80_1253 ();
 sg13g2_decap_8 FILLER_80_1260 ();
 sg13g2_decap_8 FILLER_80_1267 ();
 sg13g2_decap_8 FILLER_80_1274 ();
 sg13g2_decap_8 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1295 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_4 FILLER_80_1309 ();
 sg13g2_fill_2 FILLER_80_1313 ();
endmodule

module tt_um_crispy_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire \pcg_out[0] ;
 wire \pcg_out[1] ;
 wire \pcg_out[2] ;
 wire \pcg_out[3] ;
 wire \pcg_out[4] ;
 wire \pcg_out[5] ;
 wire \pcg_out[6] ;
 wire \pcg_out[7] ;
 wire \state[0] ;
 wire \state[10] ;
 wire \state[11] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net55;

 sg13g2_inv_1 _0731_ (.Y(_0678_),
    .A(net123));
 sg13g2_inv_1 _0732_ (.Y(_0679_),
    .A(net121));
 sg13g2_inv_1 _0733_ (.Y(_0680_),
    .A(net120));
 sg13g2_inv_1 _0734_ (.Y(_0681_),
    .A(net118));
 sg13g2_inv_1 _0735_ (.Y(_0682_),
    .A(_0008_));
 sg13g2_inv_1 _0736_ (.Y(_0683_),
    .A(\state[5] ));
 sg13g2_inv_1 _0737_ (.Y(_0684_),
    .A(net111));
 sg13g2_inv_1 _0738_ (.Y(_0685_),
    .A(_0003_));
 sg13g2_inv_1 _0739_ (.Y(_0686_),
    .A(net106));
 sg13g2_inv_2 _0740_ (.Y(_0687_),
    .A(_0004_));
 sg13g2_inv_2 _0741_ (.Y(_0688_),
    .A(net103));
 sg13g2_inv_4 _0742_ (.A(\state[15] ),
    .Y(_0689_));
 sg13g2_inv_4 _0743_ (.A(net125),
    .Y(_0690_));
 sg13g2_nand2_1 _0744_ (.Y(_0691_),
    .A(net13),
    .B(\pcg_out[4] ));
 sg13g2_xnor2_1 _0745_ (.Y(uo_out[3]),
    .A(net4),
    .B(_0691_));
 sg13g2_nand2_1 _0746_ (.Y(_0692_),
    .A(net13),
    .B(\pcg_out[5] ));
 sg13g2_nand2_1 _0747_ (.Y(_0034_),
    .A(\pcg_out[1] ),
    .B(net10));
 sg13g2_nand2_1 _0748_ (.Y(_0035_),
    .A(net9),
    .B(\pcg_out[0] ));
 sg13g2_xor2_1 _0749_ (.B(_0034_),
    .A(_0692_),
    .X(_0036_));
 sg13g2_xnor2_1 _0750_ (.Y(_0037_),
    .A(_0035_),
    .B(_0036_));
 sg13g2_nand2_1 _0751_ (.Y(_0038_),
    .A(\pcg_out[2] ),
    .B(net11));
 sg13g2_nand2_1 _0752_ (.Y(_0039_),
    .A(net14),
    .B(\pcg_out[6] ));
 sg13g2_xor2_1 _0753_ (.B(_0039_),
    .A(_0038_),
    .X(_0040_));
 sg13g2_xnor2_1 _0754_ (.Y(_0041_),
    .A(net15),
    .B(_0691_));
 sg13g2_xnor2_1 _0755_ (.Y(_0042_),
    .A(_0040_),
    .B(_0041_));
 sg13g2_nand2_1 _0756_ (.Y(_0043_),
    .A(\pcg_out[3] ),
    .B(net12));
 sg13g2_nand2_1 _0757_ (.Y(_0044_),
    .A(net14),
    .B(\pcg_out[7] ));
 sg13g2_xnor2_1 _0758_ (.Y(_0045_),
    .A(_0043_),
    .B(_0044_));
 sg13g2_xnor2_1 _0759_ (.Y(_0046_),
    .A(_0037_),
    .B(_0042_));
 sg13g2_xnor2_1 _0760_ (.Y(uio_out[7]),
    .A(_0045_),
    .B(_0046_));
 sg13g2_nand3_1 _0761_ (.B(net14),
    .C(\pcg_out[6] ),
    .A(net11),
    .Y(_0047_));
 sg13g2_xnor2_1 _0762_ (.Y(uo_out[1]),
    .A(net2),
    .B(_0047_));
 sg13g2_nand3_1 _0763_ (.B(\pcg_out[5] ),
    .C(net10),
    .A(net14),
    .Y(_0048_));
 sg13g2_xnor2_1 _0764_ (.Y(uo_out[2]),
    .A(net3),
    .B(_0048_));
 sg13g2_xnor2_1 _0765_ (.Y(uo_out[4]),
    .A(net5),
    .B(_0043_));
 sg13g2_xnor2_1 _0766_ (.Y(uo_out[5]),
    .A(net6),
    .B(_0038_));
 sg13g2_xnor2_1 _0767_ (.Y(uo_out[6]),
    .A(net7),
    .B(_0034_));
 sg13g2_xnor2_1 _0768_ (.Y(uo_out[7]),
    .A(net8),
    .B(_0035_));
 sg13g2_nand3_1 _0769_ (.B(\pcg_out[7] ),
    .C(net12),
    .A(net14),
    .Y(_0049_));
 sg13g2_xnor2_1 _0770_ (.Y(uo_out[0]),
    .A(net1),
    .B(_0049_));
 sg13g2_and2_1 _0771_ (.A(net55),
    .B(net125),
    .X(_0010_));
 sg13g2_nor2_2 _0772_ (.A(_0678_),
    .B(_0679_),
    .Y(_0050_));
 sg13g2_xor2_1 _0773_ (.B(net121),
    .A(net122),
    .X(_0051_));
 sg13g2_and2_1 _0774_ (.A(net124),
    .B(_0051_),
    .X(_0011_));
 sg13g2_nand2_2 _0775_ (.Y(_0052_),
    .A(net121),
    .B(net120));
 sg13g2_nor2_1 _0776_ (.A(net121),
    .B(net120),
    .Y(_0053_));
 sg13g2_xor2_1 _0777_ (.B(net120),
    .A(net121),
    .X(_0054_));
 sg13g2_nand2_1 _0778_ (.Y(_0055_),
    .A(net122),
    .B(_0054_));
 sg13g2_o21ai_1 _0779_ (.B1(net124),
    .Y(_0056_),
    .A1(net122),
    .A2(net120));
 sg13g2_nand2b_1 _0780_ (.Y(_0012_),
    .B(_0055_),
    .A_N(_0056_));
 sg13g2_nand3_1 _0781_ (.B(_0681_),
    .C(_0050_),
    .A(net120),
    .Y(_0057_));
 sg13g2_xor2_1 _0782_ (.B(net118),
    .A(net121),
    .X(_0058_));
 sg13g2_xnor2_1 _0783_ (.Y(_0059_),
    .A(_0680_),
    .B(_0058_));
 sg13g2_nand2_1 _0784_ (.Y(_0060_),
    .A(net122),
    .B(_0679_));
 sg13g2_a22oi_1 _0785_ (.Y(_0061_),
    .B1(_0059_),
    .B2(_0060_),
    .A2(_0058_),
    .A1(net122));
 sg13g2_nand2_1 _0786_ (.Y(_0062_),
    .A(net125),
    .B(_0057_));
 sg13g2_nor2_1 _0787_ (.A(_0061_),
    .B(_0062_),
    .Y(_0013_));
 sg13g2_nor3_2 _0788_ (.A(_0678_),
    .B(net120),
    .C(_0058_),
    .Y(_0063_));
 sg13g2_xnor2_1 _0789_ (.Y(_0064_),
    .A(net122),
    .B(_0054_));
 sg13g2_and3_1 _0790_ (.X(_0065_),
    .A(net121),
    .B(net119),
    .C(_0007_));
 sg13g2_nand3_1 _0791_ (.B(net119),
    .C(_0007_),
    .A(net121),
    .Y(_0066_));
 sg13g2_a21oi_1 _0792_ (.A1(\state[1] ),
    .A2(net119),
    .Y(_0067_),
    .B1(_0007_));
 sg13g2_nor2_1 _0793_ (.A(_0065_),
    .B(_0067_),
    .Y(_0068_));
 sg13g2_xnor2_1 _0794_ (.Y(_0069_),
    .A(_0064_),
    .B(_0068_));
 sg13g2_a22oi_1 _0795_ (.Y(_0070_),
    .B1(_0059_),
    .B2(net122),
    .A2(_0058_),
    .A1(_0682_));
 sg13g2_nand2b_1 _0796_ (.Y(_0071_),
    .B(_0070_),
    .A_N(_0069_));
 sg13g2_nor2b_1 _0797_ (.A(_0070_),
    .B_N(_0069_),
    .Y(_0072_));
 sg13g2_inv_1 _0798_ (.Y(_0073_),
    .A(_0072_));
 sg13g2_xnor2_1 _0799_ (.Y(_0074_),
    .A(_0069_),
    .B(_0070_));
 sg13g2_nand2_1 _0800_ (.Y(_0075_),
    .A(_0063_),
    .B(_0074_));
 sg13g2_inv_1 _0801_ (.Y(_0076_),
    .A(_0075_));
 sg13g2_nor2_1 _0802_ (.A(_0063_),
    .B(_0074_),
    .Y(_0077_));
 sg13g2_or2_1 _0803_ (.X(_0078_),
    .B(_0077_),
    .A(_0076_));
 sg13g2_or2_1 _0804_ (.X(_0079_),
    .B(_0078_),
    .A(_0057_));
 sg13g2_nand2_1 _0805_ (.Y(_0080_),
    .A(net125),
    .B(_0079_));
 sg13g2_a21oi_1 _0806_ (.A1(_0057_),
    .A2(_0078_),
    .Y(_0014_),
    .B1(_0080_));
 sg13g2_and2_1 _0807_ (.A(_0052_),
    .B(_0055_),
    .X(_0081_));
 sg13g2_o21ai_1 _0808_ (.B1(_0066_),
    .Y(_0082_),
    .A1(_0064_),
    .A2(_0067_));
 sg13g2_nor2b_1 _0809_ (.A(net116),
    .B_N(net117),
    .Y(_0083_));
 sg13g2_xnor2_1 _0810_ (.Y(_0084_),
    .A(net117),
    .B(net116));
 sg13g2_xor2_1 _0811_ (.B(_0084_),
    .A(_0059_),
    .X(_0085_));
 sg13g2_nand2_1 _0812_ (.Y(_0086_),
    .A(_0082_),
    .B(_0085_));
 sg13g2_xnor2_1 _0813_ (.Y(_0087_),
    .A(_0082_),
    .B(_0085_));
 sg13g2_xor2_1 _0814_ (.B(_0087_),
    .A(_0081_),
    .X(_0088_));
 sg13g2_nand2_1 _0815_ (.Y(_0089_),
    .A(_0072_),
    .B(_0088_));
 sg13g2_xnor2_1 _0816_ (.Y(_0090_),
    .A(_0072_),
    .B(_0088_));
 sg13g2_nand4_1 _0817_ (.B(_0071_),
    .C(_0073_),
    .A(_0063_),
    .Y(_0091_),
    .D(_0088_));
 sg13g2_xnor2_1 _0818_ (.Y(_0092_),
    .A(_0075_),
    .B(_0090_));
 sg13g2_nor4_2 _0819_ (.A(_0057_),
    .B(_0076_),
    .C(_0077_),
    .Y(_0093_),
    .D(_0090_));
 sg13g2_nand2b_1 _0820_ (.Y(_0094_),
    .B(net124),
    .A_N(_0093_));
 sg13g2_a21oi_1 _0821_ (.A1(_0079_),
    .A2(_0092_),
    .Y(_0015_),
    .B1(_0094_));
 sg13g2_a21oi_1 _0822_ (.A1(_0681_),
    .A2(_0052_),
    .Y(_0095_),
    .B1(_0053_));
 sg13g2_a21oi_2 _0823_ (.B1(_0083_),
    .Y(_0096_),
    .A2(_0084_),
    .A1(_0059_));
 sg13g2_and2_1 _0824_ (.A(net115),
    .B(net114),
    .X(_0097_));
 sg13g2_xor2_1 _0825_ (.B(net114),
    .A(net116),
    .X(_0098_));
 sg13g2_xnor2_1 _0826_ (.Y(_0099_),
    .A(net115),
    .B(net114));
 sg13g2_and2_1 _0827_ (.A(net118),
    .B(net117),
    .X(_0100_));
 sg13g2_xor2_1 _0828_ (.B(net117),
    .A(net118),
    .X(_0101_));
 sg13g2_xnor2_1 _0829_ (.Y(_0102_),
    .A(_0008_),
    .B(_0101_));
 sg13g2_xnor2_1 _0830_ (.Y(_0103_),
    .A(_0099_),
    .B(_0102_));
 sg13g2_nor2_1 _0831_ (.A(_0096_),
    .B(_0103_),
    .Y(_0104_));
 sg13g2_nand2_1 _0832_ (.Y(_0105_),
    .A(_0096_),
    .B(_0103_));
 sg13g2_xor2_1 _0833_ (.B(_0103_),
    .A(_0096_),
    .X(_0106_));
 sg13g2_xnor2_1 _0834_ (.Y(_0107_),
    .A(_0095_),
    .B(_0106_));
 sg13g2_o21ai_1 _0835_ (.B1(_0086_),
    .Y(_0108_),
    .A1(_0081_),
    .A2(_0087_));
 sg13g2_nand2b_1 _0836_ (.Y(_0109_),
    .B(_0108_),
    .A_N(_0107_));
 sg13g2_xor2_1 _0837_ (.B(_0108_),
    .A(_0107_),
    .X(_0110_));
 sg13g2_nand3_1 _0838_ (.B(_0091_),
    .C(_0110_),
    .A(_0089_),
    .Y(_0111_));
 sg13g2_nor2_1 _0839_ (.A(_0091_),
    .B(_0110_),
    .Y(_0112_));
 sg13g2_nor2_1 _0840_ (.A(_0089_),
    .B(_0110_),
    .Y(_0113_));
 sg13g2_a21o_1 _0841_ (.A2(_0091_),
    .A1(_0089_),
    .B1(_0110_),
    .X(_0114_));
 sg13g2_and2_1 _0842_ (.A(_0111_),
    .B(_0114_),
    .X(_0115_));
 sg13g2_nor2_1 _0843_ (.A(_0093_),
    .B(_0115_),
    .Y(_0116_));
 sg13g2_a21oi_1 _0844_ (.A1(_0093_),
    .A2(_0115_),
    .Y(_0117_),
    .B1(_0690_));
 sg13g2_nor2b_1 _0845_ (.A(_0116_),
    .B_N(_0117_),
    .Y(_0016_));
 sg13g2_a21o_1 _0846_ (.A2(_0101_),
    .A1(_0682_),
    .B1(_0100_),
    .X(_0118_));
 sg13g2_nor2_1 _0847_ (.A(_0683_),
    .B(\state[6] ),
    .Y(_0119_));
 sg13g2_a21oi_2 _0848_ (.B1(_0119_),
    .Y(_0120_),
    .A2(_0102_),
    .A1(_0099_));
 sg13g2_xnor2_1 _0849_ (.Y(_0121_),
    .A(net115),
    .B(net113));
 sg13g2_nor2_1 _0850_ (.A(_0000_),
    .B(_0121_),
    .Y(_0122_));
 sg13g2_xor2_1 _0851_ (.B(_0121_),
    .A(_0000_),
    .X(_0123_));
 sg13g2_xnor2_1 _0852_ (.Y(_0124_),
    .A(_0101_),
    .B(_0123_));
 sg13g2_nor2_1 _0853_ (.A(_0120_),
    .B(_0124_),
    .Y(_0125_));
 sg13g2_xor2_1 _0854_ (.B(_0124_),
    .A(_0120_),
    .X(_0126_));
 sg13g2_xnor2_1 _0855_ (.Y(_0127_),
    .A(_0118_),
    .B(_0126_));
 sg13g2_a21oi_1 _0856_ (.A1(_0095_),
    .A2(_0105_),
    .Y(_0128_),
    .B1(_0104_));
 sg13g2_nor2_1 _0857_ (.A(_0127_),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_xnor2_1 _0858_ (.Y(_0130_),
    .A(_0127_),
    .B(_0128_));
 sg13g2_nor2_1 _0859_ (.A(_0109_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_inv_1 _0860_ (.Y(_0132_),
    .A(_0131_));
 sg13g2_xor2_1 _0861_ (.B(_0130_),
    .A(_0109_),
    .X(_0133_));
 sg13g2_xnor2_1 _0862_ (.Y(_0134_),
    .A(_0114_),
    .B(_0133_));
 sg13g2_a21oi_1 _0863_ (.A1(_0093_),
    .A2(_0115_),
    .Y(_0135_),
    .B1(_0134_));
 sg13g2_and4_1 _0864_ (.A(_0093_),
    .B(_0111_),
    .C(_0114_),
    .D(_0133_),
    .X(_0136_));
 sg13g2_nor3_1 _0865_ (.A(_0690_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0017_));
 sg13g2_a21o_1 _0866_ (.A2(_0133_),
    .A1(_0112_),
    .B1(_0136_),
    .X(_0137_));
 sg13g2_nand2_1 _0867_ (.Y(_0138_),
    .A(_0113_),
    .B(_0133_));
 sg13g2_a21oi_1 _0868_ (.A1(_0113_),
    .A2(_0133_),
    .Y(_0139_),
    .B1(_0131_));
 sg13g2_a21oi_1 _0869_ (.A1(_0101_),
    .A2(_0123_),
    .Y(_0140_),
    .B1(_0122_));
 sg13g2_xnor2_1 _0870_ (.Y(_0141_),
    .A(net117),
    .B(_0098_));
 sg13g2_nand3_1 _0871_ (.B(net113),
    .C(_0001_),
    .A(net115),
    .Y(_0142_));
 sg13g2_a21o_1 _0872_ (.A2(net113),
    .A1(net115),
    .B1(_0001_),
    .X(_0143_));
 sg13g2_nand2_1 _0873_ (.Y(_0144_),
    .A(_0142_),
    .B(_0143_));
 sg13g2_xnor2_1 _0874_ (.Y(_0145_),
    .A(_0141_),
    .B(_0144_));
 sg13g2_nor2_1 _0875_ (.A(_0140_),
    .B(_0145_),
    .Y(_0146_));
 sg13g2_xor2_1 _0876_ (.B(_0145_),
    .A(_0140_),
    .X(_0147_));
 sg13g2_xor2_1 _0877_ (.B(_0147_),
    .A(_0100_),
    .X(_0148_));
 sg13g2_a21oi_1 _0878_ (.A1(_0118_),
    .A2(_0126_),
    .Y(_0149_),
    .B1(_0125_));
 sg13g2_nor2b_1 _0879_ (.A(_0149_),
    .B_N(_0148_),
    .Y(_0150_));
 sg13g2_inv_1 _0880_ (.Y(_0151_),
    .A(_0150_));
 sg13g2_xnor2_1 _0881_ (.Y(_0152_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_nand2_1 _0882_ (.Y(_0153_),
    .A(_0129_),
    .B(_0152_));
 sg13g2_xnor2_1 _0883_ (.Y(_0154_),
    .A(_0129_),
    .B(_0152_));
 sg13g2_xor2_1 _0884_ (.B(_0154_),
    .A(_0139_),
    .X(_0155_));
 sg13g2_xor2_1 _0885_ (.B(_0155_),
    .A(_0137_),
    .X(_0156_));
 sg13g2_nand2b_1 _0886_ (.Y(_0018_),
    .B(net124),
    .A_N(_0156_));
 sg13g2_nor2_1 _0887_ (.A(_0138_),
    .B(_0154_),
    .Y(_0157_));
 sg13g2_a21oi_2 _0888_ (.B1(_0157_),
    .Y(_0158_),
    .A2(_0155_),
    .A1(_0137_));
 sg13g2_a21oi_1 _0889_ (.A1(_0100_),
    .A2(_0147_),
    .Y(_0159_),
    .B1(_0146_));
 sg13g2_a21oi_1 _0890_ (.A1(net117),
    .A2(_0098_),
    .Y(_0160_),
    .B1(_0097_));
 sg13g2_o21ai_1 _0891_ (.B1(_0142_),
    .Y(_0161_),
    .A1(_0141_),
    .A2(_0144_));
 sg13g2_and2_1 _0892_ (.A(net112),
    .B(net111),
    .X(_0162_));
 sg13g2_xor2_1 _0893_ (.B(net111),
    .A(net112),
    .X(_0163_));
 sg13g2_and2_1 _0894_ (.A(net114),
    .B(net113),
    .X(_0164_));
 sg13g2_xor2_1 _0895_ (.B(net113),
    .A(net114),
    .X(_0165_));
 sg13g2_xnor2_1 _0896_ (.Y(_0166_),
    .A(net115),
    .B(_0165_));
 sg13g2_xor2_1 _0897_ (.B(_0166_),
    .A(_0163_),
    .X(_0167_));
 sg13g2_and2_1 _0898_ (.A(_0161_),
    .B(_0167_),
    .X(_0168_));
 sg13g2_xnor2_1 _0899_ (.Y(_0169_),
    .A(_0161_),
    .B(_0167_));
 sg13g2_nor2_1 _0900_ (.A(_0160_),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_xor2_1 _0901_ (.B(_0169_),
    .A(_0160_),
    .X(_0171_));
 sg13g2_nor2b_1 _0902_ (.A(_0159_),
    .B_N(_0171_),
    .Y(_0172_));
 sg13g2_xnor2_1 _0903_ (.Y(_0173_),
    .A(_0159_),
    .B(_0171_));
 sg13g2_xnor2_1 _0904_ (.Y(_0174_),
    .A(net123),
    .B(_0173_));
 sg13g2_or2_1 _0905_ (.X(_0175_),
    .B(_0174_),
    .A(_0151_));
 sg13g2_xnor2_1 _0906_ (.Y(_0176_),
    .A(_0151_),
    .B(_0174_));
 sg13g2_xor2_1 _0907_ (.B(_0176_),
    .A(_0153_),
    .X(_0177_));
 sg13g2_a21oi_1 _0908_ (.A1(_0131_),
    .A2(_0152_),
    .Y(_0178_),
    .B1(_0177_));
 sg13g2_nor3_1 _0909_ (.A(_0132_),
    .B(_0154_),
    .C(_0176_),
    .Y(_0179_));
 sg13g2_or3_1 _0910_ (.A(_0132_),
    .B(_0154_),
    .C(_0176_),
    .X(_0180_));
 sg13g2_o21ai_1 _0911_ (.B1(_0158_),
    .Y(_0181_),
    .A1(_0178_),
    .A2(_0179_));
 sg13g2_o21ai_1 _0912_ (.B1(net124),
    .Y(_0182_),
    .A1(_0158_),
    .A2(_0178_));
 sg13g2_nor2b_1 _0913_ (.A(_0182_),
    .B_N(_0181_),
    .Y(_0019_));
 sg13g2_o21ai_1 _0914_ (.B1(_0180_),
    .Y(_0183_),
    .A1(_0158_),
    .A2(_0178_));
 sg13g2_a21oi_1 _0915_ (.A1(net123),
    .A2(_0173_),
    .Y(_0184_),
    .B1(_0172_));
 sg13g2_a21oi_1 _0916_ (.A1(net115),
    .A2(_0165_),
    .Y(_0185_),
    .B1(_0164_));
 sg13g2_nand2_1 _0917_ (.Y(_0186_),
    .A(net112),
    .B(net109));
 sg13g2_nor2_1 _0918_ (.A(net112),
    .B(net109),
    .Y(_0187_));
 sg13g2_xor2_1 _0919_ (.B(net109),
    .A(net112),
    .X(_0188_));
 sg13g2_xnor2_1 _0920_ (.Y(_0189_),
    .A(net111),
    .B(_0188_));
 sg13g2_nor2b_1 _0921_ (.A(_0189_),
    .B_N(_0165_),
    .Y(_0190_));
 sg13g2_xnor2_1 _0922_ (.Y(_0191_),
    .A(_0165_),
    .B(_0189_));
 sg13g2_nand2_1 _0923_ (.Y(_0192_),
    .A(net112),
    .B(_0684_));
 sg13g2_o21ai_1 _0924_ (.B1(_0192_),
    .Y(_0193_),
    .A1(_0163_),
    .A2(_0166_));
 sg13g2_and2_1 _0925_ (.A(_0191_),
    .B(_0193_),
    .X(_0194_));
 sg13g2_xnor2_1 _0926_ (.Y(_0195_),
    .A(_0191_),
    .B(_0193_));
 sg13g2_nor2_1 _0927_ (.A(_0185_),
    .B(_0195_),
    .Y(_0196_));
 sg13g2_xor2_1 _0928_ (.B(_0195_),
    .A(_0185_),
    .X(_0197_));
 sg13g2_o21ai_1 _0929_ (.B1(_0197_),
    .Y(_0198_),
    .A1(_0168_),
    .A2(_0170_));
 sg13g2_nor3_1 _0930_ (.A(_0168_),
    .B(_0170_),
    .C(_0197_),
    .Y(_0199_));
 sg13g2_or3_1 _0931_ (.A(_0168_),
    .B(_0170_),
    .C(_0197_),
    .X(_0200_));
 sg13g2_and2_1 _0932_ (.A(_0198_),
    .B(_0200_),
    .X(_0201_));
 sg13g2_xnor2_1 _0933_ (.Y(_0202_),
    .A(_0002_),
    .B(_0201_));
 sg13g2_nand2b_1 _0934_ (.Y(_0203_),
    .B(_0202_),
    .A_N(_0184_));
 sg13g2_xor2_1 _0935_ (.B(_0202_),
    .A(_0184_),
    .X(_0204_));
 sg13g2_o21ai_1 _0936_ (.B1(_0175_),
    .Y(_0205_),
    .A1(_0153_),
    .A2(_0176_));
 sg13g2_xnor2_1 _0937_ (.Y(_0206_),
    .A(_0204_),
    .B(_0205_));
 sg13g2_nor2_1 _0938_ (.A(_0183_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_a21oi_1 _0939_ (.A1(_0183_),
    .A2(_0206_),
    .Y(_0208_),
    .B1(_0690_));
 sg13g2_nor2b_1 _0940_ (.A(_0207_),
    .B_N(_0208_),
    .Y(_0020_));
 sg13g2_nor3_1 _0941_ (.A(_0153_),
    .B(_0176_),
    .C(_0204_),
    .Y(_0209_));
 sg13g2_a21oi_1 _0942_ (.A1(_0183_),
    .A2(_0206_),
    .Y(_0210_),
    .B1(_0209_));
 sg13g2_nor3_1 _0943_ (.A(_0151_),
    .B(_0174_),
    .C(_0204_),
    .Y(_0211_));
 sg13g2_a21oi_1 _0944_ (.A1(_0685_),
    .A2(_0188_),
    .Y(_0212_),
    .B1(_0190_));
 sg13g2_xnor2_1 _0945_ (.Y(_0213_),
    .A(net113),
    .B(_0163_));
 sg13g2_nand2_1 _0946_ (.Y(_0214_),
    .A(net110),
    .B(\state[11] ));
 sg13g2_xor2_1 _0947_ (.B(_0186_),
    .A(net108),
    .X(_0215_));
 sg13g2_nand2b_1 _0948_ (.Y(_0216_),
    .B(_0215_),
    .A_N(_0213_));
 sg13g2_xor2_1 _0949_ (.B(_0215_),
    .A(_0213_),
    .X(_0217_));
 sg13g2_nor2_1 _0950_ (.A(_0212_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_xor2_1 _0951_ (.B(_0217_),
    .A(_0212_),
    .X(_0219_));
 sg13g2_xor2_1 _0952_ (.B(_0219_),
    .A(_0164_),
    .X(_0220_));
 sg13g2_nor3_1 _0953_ (.A(_0194_),
    .B(_0196_),
    .C(_0220_),
    .Y(_0221_));
 sg13g2_o21ai_1 _0954_ (.B1(_0220_),
    .Y(_0222_),
    .A1(_0194_),
    .A2(_0196_));
 sg13g2_nor2b_1 _0955_ (.A(_0221_),
    .B_N(_0222_),
    .Y(_0223_));
 sg13g2_xnor2_1 _0956_ (.Y(_0224_),
    .A(_0008_),
    .B(_0223_));
 sg13g2_o21ai_1 _0957_ (.B1(_0198_),
    .Y(_0225_),
    .A1(_0679_),
    .A2(_0199_));
 sg13g2_xnor2_1 _0958_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_nor2_1 _0959_ (.A(_0203_),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_xor2_1 _0960_ (.B(_0226_),
    .A(_0203_),
    .X(_0228_));
 sg13g2_nand2_1 _0961_ (.Y(_0229_),
    .A(_0211_),
    .B(_0228_));
 sg13g2_xnor2_1 _0962_ (.Y(_0230_),
    .A(_0211_),
    .B(_0228_));
 sg13g2_o21ai_1 _0963_ (.B1(net124),
    .Y(_0231_),
    .A1(_0210_),
    .A2(_0230_));
 sg13g2_a21oi_1 _0964_ (.A1(_0210_),
    .A2(_0230_),
    .Y(_0021_),
    .B1(_0231_));
 sg13g2_o21ai_1 _0965_ (.B1(_0229_),
    .Y(_0232_),
    .A1(_0210_),
    .A2(_0230_));
 sg13g2_nand2_2 _0966_ (.Y(_0233_),
    .A(net122),
    .B(net118));
 sg13g2_xor2_1 _0967_ (.B(net118),
    .A(net123),
    .X(_0234_));
 sg13g2_a21oi_1 _0968_ (.A1(_0164_),
    .A2(_0219_),
    .Y(_0235_),
    .B1(_0218_));
 sg13g2_a21oi_1 _0969_ (.A1(net113),
    .A2(_0163_),
    .Y(_0236_),
    .B1(_0162_));
 sg13g2_xnor2_1 _0970_ (.Y(_0237_),
    .A(net108),
    .B(net106));
 sg13g2_nor2b_1 _0971_ (.A(_0189_),
    .B_N(_0237_),
    .Y(_0238_));
 sg13g2_xnor2_1 _0972_ (.Y(_0239_),
    .A(_0189_),
    .B(_0237_));
 sg13g2_o21ai_1 _0973_ (.B1(_0216_),
    .Y(_0240_),
    .A1(_0687_),
    .A2(_0186_));
 sg13g2_xor2_1 _0974_ (.B(_0240_),
    .A(_0239_),
    .X(_0241_));
 sg13g2_nor2b_1 _0975_ (.A(_0236_),
    .B_N(_0241_),
    .Y(_0242_));
 sg13g2_xnor2_1 _0976_ (.Y(_0243_),
    .A(_0236_),
    .B(_0241_));
 sg13g2_nor2b_1 _0977_ (.A(_0235_),
    .B_N(_0243_),
    .Y(_0244_));
 sg13g2_xnor2_1 _0978_ (.Y(_0245_),
    .A(_0235_),
    .B(_0243_));
 sg13g2_xnor2_1 _0979_ (.Y(_0246_),
    .A(_0234_),
    .B(_0245_));
 sg13g2_a21oi_1 _0980_ (.A1(_0680_),
    .A2(_0222_),
    .Y(_0247_),
    .B1(_0221_));
 sg13g2_nand2b_1 _0981_ (.Y(_0248_),
    .B(_0247_),
    .A_N(_0246_));
 sg13g2_xnor2_1 _0982_ (.Y(_0249_),
    .A(_0246_),
    .B(_0247_));
 sg13g2_a21oi_1 _0983_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0250_),
    .B1(_0227_));
 sg13g2_xnor2_1 _0984_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_xnor2_1 _0985_ (.Y(_0252_),
    .A(_0232_),
    .B(_0251_));
 sg13g2_nand2_1 _0986_ (.Y(_0022_),
    .A(net124),
    .B(_0252_));
 sg13g2_a22oi_1 _0987_ (.Y(_0253_),
    .B1(_0251_),
    .B2(_0232_),
    .A2(_0249_),
    .A1(_0227_));
 sg13g2_a21o_1 _0988_ (.A2(_0240_),
    .A1(_0239_),
    .B1(_0242_),
    .X(_0254_));
 sg13g2_a21oi_1 _0989_ (.A1(_0684_),
    .A2(_0186_),
    .Y(_0255_),
    .B1(_0187_));
 sg13g2_a21oi_1 _0990_ (.A1(net108),
    .A2(_0686_),
    .Y(_0256_),
    .B1(_0238_));
 sg13g2_or2_1 _0991_ (.X(_0257_),
    .B(net104),
    .A(net106));
 sg13g2_xor2_1 _0992_ (.B(net103),
    .A(net106),
    .X(_0258_));
 sg13g2_nor2_1 _0993_ (.A(net110),
    .B(\state[11] ),
    .Y(_0259_));
 sg13g2_xor2_1 _0994_ (.B(net108),
    .A(net110),
    .X(_0260_));
 sg13g2_inv_1 _0995_ (.Y(_0261_),
    .A(_0260_));
 sg13g2_xnor2_1 _0996_ (.Y(_0262_),
    .A(net111),
    .B(_0260_));
 sg13g2_xnor2_1 _0997_ (.Y(_0263_),
    .A(_0258_),
    .B(_0262_));
 sg13g2_nor2_1 _0998_ (.A(_0256_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_nand2_1 _0999_ (.Y(_0265_),
    .A(_0256_),
    .B(_0263_));
 sg13g2_nand2b_1 _1000_ (.Y(_0266_),
    .B(_0265_),
    .A_N(_0264_));
 sg13g2_xor2_1 _1001_ (.B(_0266_),
    .A(_0255_),
    .X(_0267_));
 sg13g2_inv_1 _1002_ (.Y(_0268_),
    .A(_0267_));
 sg13g2_xnor2_1 _1003_ (.Y(_0269_),
    .A(_0254_),
    .B(_0268_));
 sg13g2_nand2_1 _1004_ (.Y(_0270_),
    .A(\state[4] ),
    .B(_0051_));
 sg13g2_xnor2_1 _1005_ (.Y(_0271_),
    .A(net117),
    .B(_0051_));
 sg13g2_or2_1 _1006_ (.X(_0272_),
    .B(_0271_),
    .A(_0233_));
 sg13g2_xnor2_1 _1007_ (.Y(_0273_),
    .A(_0233_),
    .B(_0271_));
 sg13g2_nor2_1 _1008_ (.A(_0269_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_xor2_1 _1009_ (.B(_0273_),
    .A(_0269_),
    .X(_0275_));
 sg13g2_a21o_1 _1010_ (.A2(_0245_),
    .A1(_0234_),
    .B1(_0244_),
    .X(_0276_));
 sg13g2_nand2_1 _1011_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_xor2_1 _1012_ (.B(_0276_),
    .A(_0275_),
    .X(_0278_));
 sg13g2_and3_1 _1013_ (.X(_0279_),
    .A(_0224_),
    .B(_0225_),
    .C(_0249_));
 sg13g2_inv_1 _1014_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nand2_1 _1015_ (.Y(_0281_),
    .A(_0248_),
    .B(_0280_));
 sg13g2_xnor2_1 _1016_ (.Y(_0282_),
    .A(_0278_),
    .B(_0281_));
 sg13g2_or2_1 _1017_ (.X(_0283_),
    .B(_0282_),
    .A(_0253_));
 sg13g2_a21oi_1 _1018_ (.A1(_0253_),
    .A2(_0282_),
    .Y(_0284_),
    .B1(_0690_));
 sg13g2_and2_1 _1019_ (.A(_0283_),
    .B(_0284_),
    .X(_0023_));
 sg13g2_nor2b_1 _1020_ (.A(_0248_),
    .B_N(_0278_),
    .Y(_0285_));
 sg13g2_a21oi_1 _1021_ (.A1(_0254_),
    .A2(_0268_),
    .Y(_0286_),
    .B1(_0274_));
 sg13g2_a21oi_1 _1022_ (.A1(_0255_),
    .A2(_0265_),
    .Y(_0287_),
    .B1(_0264_));
 sg13g2_nand2_1 _1023_ (.Y(_0288_),
    .A(net106),
    .B(_0688_));
 sg13g2_o21ai_1 _1024_ (.B1(_0288_),
    .Y(_0289_),
    .A1(_0258_),
    .A2(_0262_));
 sg13g2_nand2_1 _1025_ (.Y(_0290_),
    .A(net107),
    .B(net99));
 sg13g2_nor2_1 _1026_ (.A(net107),
    .B(net100),
    .Y(_0291_));
 sg13g2_xor2_1 _1027_ (.B(net99),
    .A(net106),
    .X(_0292_));
 sg13g2_xnor2_1 _1028_ (.Y(_0293_),
    .A(net104),
    .B(_0292_));
 sg13g2_nor2_1 _1029_ (.A(_0261_),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_xnor2_1 _1030_ (.Y(_0295_),
    .A(_0260_),
    .B(_0293_));
 sg13g2_and2_1 _1031_ (.A(_0289_),
    .B(_0295_),
    .X(_0296_));
 sg13g2_xor2_1 _1032_ (.B(_0295_),
    .A(_0289_),
    .X(_0297_));
 sg13g2_a21oi_1 _1033_ (.A1(_0003_),
    .A2(_0214_),
    .Y(_0298_),
    .B1(_0259_));
 sg13g2_xnor2_1 _1034_ (.Y(_0299_),
    .A(_0297_),
    .B(_0298_));
 sg13g2_nor2_1 _1035_ (.A(_0287_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_xor2_1 _1036_ (.B(_0299_),
    .A(_0287_),
    .X(_0301_));
 sg13g2_xnor2_1 _1037_ (.Y(_0302_),
    .A(net115),
    .B(_0054_));
 sg13g2_nor2_1 _1038_ (.A(_0270_),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_xor2_1 _1039_ (.B(_0302_),
    .A(_0270_),
    .X(_0304_));
 sg13g2_xnor2_1 _1040_ (.Y(_0305_),
    .A(_0301_),
    .B(_0304_));
 sg13g2_or2_1 _1041_ (.X(_0306_),
    .B(_0305_),
    .A(_0286_));
 sg13g2_xnor2_1 _1042_ (.Y(_0307_),
    .A(_0286_),
    .B(_0305_));
 sg13g2_xnor2_1 _1043_ (.Y(_0308_),
    .A(_0272_),
    .B(_0307_));
 sg13g2_nor2_1 _1044_ (.A(_0277_),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_xor2_1 _1045_ (.B(_0308_),
    .A(_0277_),
    .X(_0310_));
 sg13g2_xor2_1 _1046_ (.B(_0310_),
    .A(_0050_),
    .X(_0311_));
 sg13g2_nand2_1 _1047_ (.Y(_0312_),
    .A(_0285_),
    .B(_0311_));
 sg13g2_xnor2_1 _1048_ (.Y(_0313_),
    .A(_0285_),
    .B(_0311_));
 sg13g2_nand2_1 _1049_ (.Y(_0314_),
    .A(_0278_),
    .B(_0279_));
 sg13g2_and2_1 _1050_ (.A(_0283_),
    .B(_0314_),
    .X(_0315_));
 sg13g2_or2_1 _1051_ (.X(_0316_),
    .B(_0315_),
    .A(_0313_));
 sg13g2_nand2_1 _1052_ (.Y(_0317_),
    .A(net124),
    .B(_0316_));
 sg13g2_a21oi_1 _1053_ (.A1(_0313_),
    .A2(_0315_),
    .Y(_0024_),
    .B1(_0317_));
 sg13g2_a21oi_1 _1054_ (.A1(_0050_),
    .A2(_0310_),
    .Y(_0318_),
    .B1(_0309_));
 sg13g2_o21ai_1 _1055_ (.B1(_0306_),
    .Y(_0319_),
    .A1(_0272_),
    .A2(_0307_));
 sg13g2_a21oi_1 _1056_ (.A1(_0301_),
    .A2(_0304_),
    .Y(_0320_),
    .B1(_0300_));
 sg13g2_xor2_1 _1057_ (.B(_0214_),
    .A(net114),
    .X(_0321_));
 sg13g2_xnor2_1 _1058_ (.Y(_0322_),
    .A(_0689_),
    .B(_0290_));
 sg13g2_xnor2_1 _1059_ (.Y(_0323_),
    .A(_0321_),
    .B(_0322_));
 sg13g2_xnor2_1 _1060_ (.Y(_0324_),
    .A(_0688_),
    .B(_0237_));
 sg13g2_xnor2_1 _1061_ (.Y(_0325_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_xor2_1 _1062_ (.B(net119),
    .A(net120),
    .X(_0326_));
 sg13g2_a21oi_2 _1063_ (.B1(_0303_),
    .Y(_0327_),
    .A2(_0054_),
    .A1(\state[5] ));
 sg13g2_a21oi_1 _1064_ (.A1(net104),
    .A2(_0292_),
    .Y(_0328_),
    .B1(_0294_));
 sg13g2_xnor2_1 _1065_ (.Y(_0329_),
    .A(_0326_),
    .B(_0328_));
 sg13g2_xnor2_1 _1066_ (.Y(_0330_),
    .A(_0325_),
    .B(_0327_));
 sg13g2_xnor2_1 _1067_ (.Y(_0331_),
    .A(_0329_),
    .B(_0330_));
 sg13g2_a21oi_1 _1068_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0332_),
    .B1(_0296_));
 sg13g2_xor2_1 _1069_ (.B(_0332_),
    .A(_0052_),
    .X(_0333_));
 sg13g2_xnor2_1 _1070_ (.Y(_0334_),
    .A(_0331_),
    .B(_0333_));
 sg13g2_xnor2_1 _1071_ (.Y(_0335_),
    .A(_0320_),
    .B(_0334_));
 sg13g2_xnor2_1 _1072_ (.Y(_0336_),
    .A(_0319_),
    .B(_0335_));
 sg13g2_xnor2_1 _1073_ (.Y(_0337_),
    .A(_0318_),
    .B(_0336_));
 sg13g2_a21oi_1 _1074_ (.A1(_0312_),
    .A2(_0316_),
    .Y(_0338_),
    .B1(_0337_));
 sg13g2_and3_1 _1075_ (.X(_0339_),
    .A(_0312_),
    .B(_0316_),
    .C(_0337_));
 sg13g2_nor3_1 _1076_ (.A(_0690_),
    .B(_0338_),
    .C(_0339_),
    .Y(_0025_));
 sg13g2_mux2_1 _1077_ (.A0(\state[7] ),
    .A1(\state[8] ),
    .S(net101),
    .X(_0340_));
 sg13g2_mux2_1 _1078_ (.A0(\state[9] ),
    .A1(net109),
    .S(net101),
    .X(_0341_));
 sg13g2_mux4_1 _1079_ (.S0(net101),
    .A0(\state[7] ),
    .A1(\state[8] ),
    .A2(\state[9] ),
    .A3(net109),
    .S1(net97),
    .X(_0342_));
 sg13g2_nor2_1 _1080_ (.A(net98),
    .B(net96),
    .Y(_0343_));
 sg13g2_nor2_1 _1081_ (.A(net117),
    .B(_0688_),
    .Y(_0344_));
 sg13g2_o21ai_1 _1082_ (.B1(_0343_),
    .Y(_0345_),
    .A1(net118),
    .A2(net102));
 sg13g2_nor2b_1 _1083_ (.A(net96),
    .B_N(net97),
    .Y(_0346_));
 sg13g2_mux2_1 _1084_ (.A0(net116),
    .A1(\state[6] ),
    .S(net101),
    .X(_0347_));
 sg13g2_a22oi_1 _1085_ (.Y(_0348_),
    .B1(_0346_),
    .B2(_0347_),
    .A2(_0342_),
    .A1(net96));
 sg13g2_o21ai_1 _1086_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_xor2_1 _1087_ (.B(_0349_),
    .A(_0009_),
    .X(_0350_));
 sg13g2_mux2_1 _1088_ (.A0(net112),
    .A1(net111),
    .S(net101),
    .X(_0351_));
 sg13g2_mux2_1 _1089_ (.A0(net109),
    .A1(net108),
    .S(net101),
    .X(_0352_));
 sg13g2_mux4_1 _1090_ (.S0(net101),
    .A0(net112),
    .A1(net111),
    .A2(net110),
    .A3(net108),
    .S1(net97),
    .X(_0353_));
 sg13g2_mux2_1 _1091_ (.A0(net114),
    .A1(\state[7] ),
    .S(net102),
    .X(_0354_));
 sg13g2_mux2_1 _1092_ (.A0(\state[4] ),
    .A1(net116),
    .S(net101),
    .X(_0355_));
 sg13g2_mux4_1 _1093_ (.S0(net97),
    .A0(_0351_),
    .A1(_0352_),
    .A2(_0355_),
    .A3(_0354_),
    .S1(_0689_),
    .X(_0356_));
 sg13g2_xnor2_1 _1094_ (.Y(_0357_),
    .A(\state[1] ),
    .B(_0356_));
 sg13g2_nor2_2 _1095_ (.A(_0350_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_nor2_1 _1096_ (.A(\state[15] ),
    .B(_0353_),
    .Y(_0359_));
 sg13g2_or2_1 _1097_ (.X(_0360_),
    .B(_0353_),
    .A(net96));
 sg13g2_nor2b_2 _1098_ (.A(net105),
    .B_N(\state[15] ),
    .Y(_0361_));
 sg13g2_and2_1 _1099_ (.A(_0291_),
    .B(_0361_),
    .X(_0362_));
 sg13g2_nand2_1 _1100_ (.Y(_0363_),
    .A(_0291_),
    .B(_0361_));
 sg13g2_a21oi_2 _1101_ (.B1(_0683_),
    .Y(_0364_),
    .A2(_0363_),
    .A1(_0360_));
 sg13g2_o21ai_1 _1102_ (.B1(net116),
    .Y(_0365_),
    .A1(_0359_),
    .A2(_0362_));
 sg13g2_nor3_2 _1103_ (.A(net116),
    .B(_0359_),
    .C(_0362_),
    .Y(_0366_));
 sg13g2_nand3_1 _1104_ (.B(_0360_),
    .C(_0363_),
    .A(_0683_),
    .Y(_0367_));
 sg13g2_nor2_2 _1105_ (.A(_0364_),
    .B(_0366_),
    .Y(_0368_));
 sg13g2_xnor2_1 _1106_ (.Y(_0369_),
    .A(_0002_),
    .B(_0356_));
 sg13g2_mux2_1 _1107_ (.A0(net108),
    .A1(net106),
    .S(net102),
    .X(_0370_));
 sg13g2_mux4_1 _1108_ (.S0(net103),
    .A0(net111),
    .A1(net109),
    .A2(net108),
    .A3(net106),
    .S1(net99),
    .X(_0371_));
 sg13g2_mux4_1 _1109_ (.S0(_0689_),
    .A0(_0341_),
    .A1(_0347_),
    .A2(_0370_),
    .A3(_0340_),
    .S1(net98),
    .X(_0372_));
 sg13g2_xnor2_1 _1110_ (.Y(_0373_),
    .A(\state[2] ),
    .B(_0372_));
 sg13g2_xor2_1 _1111_ (.B(_0373_),
    .A(_0369_),
    .X(_0374_));
 sg13g2_nor2_1 _1112_ (.A(_0368_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_xnor2_1 _1113_ (.Y(_0376_),
    .A(_0368_),
    .B(_0374_));
 sg13g2_xnor2_1 _1114_ (.Y(_0377_),
    .A(_0358_),
    .B(_0376_));
 sg13g2_mux2_1 _1115_ (.A0(_0352_),
    .A1(_0257_),
    .S(net97),
    .X(_0378_));
 sg13g2_mux4_1 _1116_ (.S0(net96),
    .A0(_0354_),
    .A1(_0352_),
    .A2(_0351_),
    .A3(_0257_),
    .S1(net97),
    .X(_0379_));
 sg13g2_xnor2_1 _1117_ (.Y(_0380_),
    .A(net118),
    .B(_0379_));
 sg13g2_nor2_1 _1118_ (.A(_0350_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_inv_1 _1119_ (.Y(_0382_),
    .A(_0381_));
 sg13g2_xnor2_1 _1120_ (.Y(_0383_),
    .A(net95),
    .B(_0357_));
 sg13g2_mux2_1 _1121_ (.A0(_0370_),
    .A1(net104),
    .S(net97),
    .X(_0384_));
 sg13g2_mux4_1 _1122_ (.S0(net97),
    .A0(_0340_),
    .A1(_0341_),
    .A2(_0370_),
    .A3(net104),
    .S1(net96),
    .X(_0385_));
 sg13g2_xnor2_1 _1123_ (.Y(_0386_),
    .A(_0007_),
    .B(_0385_));
 sg13g2_xor2_1 _1124_ (.B(_0385_),
    .A(_0007_),
    .X(_0387_));
 sg13g2_nand2b_2 _1125_ (.Y(_0388_),
    .B(_0386_),
    .A_N(_0383_));
 sg13g2_xnor2_1 _1126_ (.Y(_0389_),
    .A(_0383_),
    .B(_0386_));
 sg13g2_xnor2_1 _1127_ (.Y(_0390_),
    .A(_0008_),
    .B(_0372_));
 sg13g2_nand2_2 _1128_ (.Y(_0391_),
    .A(_0369_),
    .B(_0390_));
 sg13g2_nor2_1 _1129_ (.A(net95),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_nand2b_2 _1130_ (.Y(_0393_),
    .B(_0390_),
    .A_N(_0380_));
 sg13g2_xnor2_1 _1131_ (.Y(_0394_),
    .A(_0380_),
    .B(_0390_));
 sg13g2_a22oi_1 _1132_ (.Y(_0395_),
    .B1(_0371_),
    .B2(_0689_),
    .A2(_0361_),
    .A1(net98));
 sg13g2_xor2_1 _1133_ (.B(_0395_),
    .A(net114),
    .X(_0396_));
 sg13g2_xnor2_1 _1134_ (.Y(_0397_),
    .A(\state[6] ),
    .B(_0395_));
 sg13g2_nand2_1 _1135_ (.Y(_0398_),
    .A(_0394_),
    .B(_0397_));
 sg13g2_xnor2_1 _1136_ (.Y(_0399_),
    .A(_0394_),
    .B(_0396_));
 sg13g2_and2_1 _1137_ (.A(_0375_),
    .B(_0399_),
    .X(_0400_));
 sg13g2_xor2_1 _1138_ (.B(_0391_),
    .A(net95),
    .X(_0401_));
 sg13g2_or2_1 _1139_ (.X(_0402_),
    .B(_0399_),
    .A(_0375_));
 sg13g2_nand2b_1 _1140_ (.Y(_0403_),
    .B(_0402_),
    .A_N(_0400_));
 sg13g2_a21o_1 _1141_ (.A2(_0402_),
    .A1(_0401_),
    .B1(_0400_),
    .X(_0404_));
 sg13g2_nor2_1 _1142_ (.A(_0383_),
    .B(_0393_),
    .Y(_0405_));
 sg13g2_xor2_1 _1143_ (.B(_0393_),
    .A(_0383_),
    .X(_0406_));
 sg13g2_nor2_1 _1144_ (.A(_0380_),
    .B(_0387_),
    .Y(_0407_));
 sg13g2_inv_1 _1145_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_xnor2_1 _1146_ (.Y(_0409_),
    .A(_0380_),
    .B(_0387_));
 sg13g2_o21ai_1 _1147_ (.B1(net96),
    .Y(_0410_),
    .A1(_0688_),
    .A2(net98));
 sg13g2_o21ai_1 _1148_ (.B1(_0410_),
    .Y(_0411_),
    .A1(net96),
    .A2(_0378_));
 sg13g2_xor2_1 _1149_ (.B(_0411_),
    .A(net113),
    .X(_0412_));
 sg13g2_nor2_1 _1150_ (.A(_0409_),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_xnor2_1 _1151_ (.Y(_0414_),
    .A(_0409_),
    .B(_0412_));
 sg13g2_nor2_1 _1152_ (.A(_0398_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_xor2_1 _1153_ (.B(_0414_),
    .A(_0398_),
    .X(_0416_));
 sg13g2_xnor2_1 _1154_ (.Y(_0417_),
    .A(_0406_),
    .B(_0416_));
 sg13g2_nor2b_1 _1155_ (.A(_0417_),
    .B_N(_0404_),
    .Y(_0418_));
 sg13g2_xnor2_1 _1156_ (.Y(_0419_),
    .A(_0404_),
    .B(_0417_));
 sg13g2_xor2_1 _1157_ (.B(_0403_),
    .A(_0401_),
    .X(_0420_));
 sg13g2_xnor2_1 _1158_ (.Y(_0421_),
    .A(_0392_),
    .B(_0419_));
 sg13g2_nor2_1 _1159_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_nand4_1 _1160_ (.B(_0381_),
    .C(_0389_),
    .A(_0377_),
    .Y(_0423_),
    .D(_0422_));
 sg13g2_nor2b_1 _1161_ (.A(_0358_),
    .B_N(_0388_),
    .Y(_0424_));
 sg13g2_nor4_2 _1162_ (.A(_0376_),
    .B(_0420_),
    .C(_0421_),
    .Y(_0425_),
    .D(_0424_));
 sg13g2_a21oi_1 _1163_ (.A1(_0406_),
    .A2(_0416_),
    .Y(_0426_),
    .B1(_0415_));
 sg13g2_a21oi_2 _1164_ (.B1(_0387_),
    .Y(_0427_),
    .A2(_0367_),
    .A1(_0365_));
 sg13g2_nor3_2 _1165_ (.A(_0364_),
    .B(_0366_),
    .C(_0386_),
    .Y(_0428_));
 sg13g2_nor2_1 _1166_ (.A(_0427_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_a22oi_1 _1167_ (.Y(_0430_),
    .B1(_0384_),
    .B2(_0689_),
    .A2(_0361_),
    .A1(_0005_));
 sg13g2_xnor2_1 _1168_ (.Y(_0431_),
    .A(_0001_),
    .B(_0430_));
 sg13g2_or3_2 _1169_ (.A(_0427_),
    .B(_0428_),
    .C(_0431_),
    .X(_0432_));
 sg13g2_o21ai_1 _1170_ (.B1(_0431_),
    .Y(_0433_),
    .A1(_0427_),
    .A2(_0428_));
 sg13g2_nand3_1 _1171_ (.B(_0432_),
    .C(_0433_),
    .A(_0413_),
    .Y(_0434_));
 sg13g2_a21oi_1 _1172_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0435_),
    .B1(_0413_));
 sg13g2_a21o_1 _1173_ (.A2(_0433_),
    .A1(_0432_),
    .B1(_0413_),
    .X(_0436_));
 sg13g2_nor2_1 _1174_ (.A(_0374_),
    .B(_0408_),
    .Y(_0437_));
 sg13g2_xnor2_1 _1175_ (.Y(_0438_),
    .A(_0374_),
    .B(_0407_));
 sg13g2_xor2_1 _1176_ (.B(_0438_),
    .A(_0358_),
    .X(_0439_));
 sg13g2_xnor2_1 _1177_ (.Y(_0440_),
    .A(_0358_),
    .B(_0438_));
 sg13g2_and3_1 _1178_ (.X(_0441_),
    .A(_0434_),
    .B(_0436_),
    .C(_0439_));
 sg13g2_a21oi_1 _1179_ (.A1(_0434_),
    .A2(_0436_),
    .Y(_0442_),
    .B1(_0439_));
 sg13g2_nor3_1 _1180_ (.A(_0426_),
    .B(_0441_),
    .C(_0442_),
    .Y(_0443_));
 sg13g2_o21ai_1 _1181_ (.B1(_0426_),
    .Y(_0444_),
    .A1(_0441_),
    .A2(_0442_));
 sg13g2_nand2b_1 _1182_ (.Y(_0445_),
    .B(_0444_),
    .A_N(_0443_));
 sg13g2_xnor2_1 _1183_ (.Y(_0446_),
    .A(_0405_),
    .B(_0445_));
 sg13g2_a21oi_1 _1184_ (.A1(_0392_),
    .A2(_0419_),
    .Y(_0447_),
    .B1(_0418_));
 sg13g2_nor2b_1 _1185_ (.A(_0447_),
    .B_N(_0446_),
    .Y(_0448_));
 sg13g2_xnor2_1 _1186_ (.Y(_0449_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_xnor2_1 _1187_ (.Y(_0450_),
    .A(_0425_),
    .B(_0449_));
 sg13g2_and2_1 _1188_ (.A(_0423_),
    .B(_0450_),
    .X(_0451_));
 sg13g2_nor2_2 _1189_ (.A(_0423_),
    .B(_0450_),
    .Y(_0452_));
 sg13g2_nor3_1 _1190_ (.A(_0690_),
    .B(_0451_),
    .C(_0452_),
    .Y(_0026_));
 sg13g2_o21ai_1 _1191_ (.B1(net95),
    .Y(_0453_),
    .A1(_0374_),
    .A2(_0408_));
 sg13g2_a21oi_1 _1192_ (.A1(_0358_),
    .A2(_0438_),
    .Y(_0454_),
    .B1(_0437_));
 sg13g2_or2_2 _1193_ (.X(_0455_),
    .B(_0454_),
    .A(net95));
 sg13g2_o21ai_1 _1194_ (.B1(_0434_),
    .Y(_0456_),
    .A1(_0435_),
    .A2(_0440_));
 sg13g2_nand2_1 _1195_ (.Y(_0457_),
    .A(_0394_),
    .B(_0427_));
 sg13g2_xnor2_1 _1196_ (.Y(_0458_),
    .A(_0394_),
    .B(_0427_));
 sg13g2_or2_1 _1197_ (.X(_0459_),
    .B(_0458_),
    .A(_0391_));
 sg13g2_xor2_1 _1198_ (.B(_0458_),
    .A(_0391_),
    .X(_0460_));
 sg13g2_nor2_1 _1199_ (.A(_0368_),
    .B(_0396_),
    .Y(_0461_));
 sg13g2_o21ai_1 _1200_ (.B1(_0397_),
    .Y(_0462_),
    .A1(_0364_),
    .A2(_0366_));
 sg13g2_nand3_1 _1201_ (.B(_0367_),
    .C(_0396_),
    .A(_0365_),
    .Y(_0463_));
 sg13g2_nand2_1 _1202_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_and2_1 _1203_ (.A(_0688_),
    .B(_0346_),
    .X(_0465_));
 sg13g2_a21o_1 _1204_ (.A2(_0343_),
    .A1(_0257_),
    .B1(_0465_),
    .X(_0466_));
 sg13g2_xnor2_1 _1205_ (.Y(_0467_),
    .A(_0003_),
    .B(_0466_));
 sg13g2_xnor2_1 _1206_ (.Y(_0468_),
    .A(_0685_),
    .B(_0466_));
 sg13g2_and3_1 _1207_ (.X(_0469_),
    .A(_0462_),
    .B(_0463_),
    .C(_0467_));
 sg13g2_a21oi_1 _1208_ (.A1(_0462_),
    .A2(_0463_),
    .Y(_0470_),
    .B1(_0467_));
 sg13g2_or3_1 _1209_ (.A(_0432_),
    .B(_0469_),
    .C(_0470_),
    .X(_0471_));
 sg13g2_o21ai_1 _1210_ (.B1(_0432_),
    .Y(_0472_),
    .A1(_0469_),
    .A2(_0470_));
 sg13g2_nand3_1 _1211_ (.B(_0471_),
    .C(_0472_),
    .A(_0460_),
    .Y(_0473_));
 sg13g2_a21o_1 _1212_ (.A2(_0472_),
    .A1(_0471_),
    .B1(_0460_),
    .X(_0474_));
 sg13g2_nand3_1 _1213_ (.B(_0473_),
    .C(_0474_),
    .A(_0456_),
    .Y(_0475_));
 sg13g2_a21o_1 _1214_ (.A2(_0474_),
    .A1(_0473_),
    .B1(_0456_),
    .X(_0476_));
 sg13g2_and4_1 _1215_ (.A(_0453_),
    .B(_0455_),
    .C(_0475_),
    .D(_0476_),
    .X(_0477_));
 sg13g2_nand4_1 _1216_ (.B(_0455_),
    .C(_0475_),
    .A(_0453_),
    .Y(_0478_),
    .D(_0476_));
 sg13g2_a22oi_1 _1217_ (.Y(_0479_),
    .B1(_0475_),
    .B2(_0476_),
    .A2(_0455_),
    .A1(_0453_));
 sg13g2_a21oi_1 _1218_ (.A1(_0405_),
    .A2(_0444_),
    .Y(_0480_),
    .B1(_0443_));
 sg13g2_o21ai_1 _1219_ (.B1(_0480_),
    .Y(_0481_),
    .A1(_0477_),
    .A2(_0479_));
 sg13g2_or3_1 _1220_ (.A(_0477_),
    .B(_0479_),
    .C(_0480_),
    .X(_0482_));
 sg13g2_and2_1 _1221_ (.A(_0481_),
    .B(_0482_),
    .X(_0483_));
 sg13g2_nand3_1 _1222_ (.B(_0449_),
    .C(_0483_),
    .A(_0425_),
    .Y(_0484_));
 sg13g2_inv_1 _1223_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_a221oi_1 _1224_ (.B2(_0482_),
    .C1(_0448_),
    .B1(_0481_),
    .A1(_0425_),
    .Y(_0486_),
    .A2(_0449_));
 sg13g2_and2_1 _1225_ (.A(_0448_),
    .B(_0483_),
    .X(_0487_));
 sg13g2_nor2_1 _1226_ (.A(_0486_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_and2_1 _1227_ (.A(_0484_),
    .B(_0488_),
    .X(_0489_));
 sg13g2_o21ai_1 _1228_ (.B1(net126),
    .Y(_0490_),
    .A1(_0452_),
    .A2(_0489_));
 sg13g2_a21oi_1 _1229_ (.A1(_0452_),
    .A2(_0489_),
    .Y(_0027_),
    .B1(_0490_));
 sg13g2_nand2_1 _1230_ (.Y(_0491_),
    .A(_0475_),
    .B(_0478_));
 sg13g2_a21o_1 _1231_ (.A2(_0459_),
    .A1(_0457_),
    .B1(_0357_),
    .X(_0492_));
 sg13g2_nand3_1 _1232_ (.B(_0457_),
    .C(_0459_),
    .A(_0357_),
    .Y(_0493_));
 sg13g2_nand2_1 _1233_ (.Y(_0494_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_nand2_1 _1234_ (.Y(_0495_),
    .A(_0471_),
    .B(_0473_));
 sg13g2_or2_1 _1235_ (.X(_0496_),
    .B(_0462_),
    .A(_0409_));
 sg13g2_xnor2_1 _1236_ (.Y(_0497_),
    .A(_0409_),
    .B(_0462_));
 sg13g2_or2_1 _1237_ (.X(_0498_),
    .B(_0497_),
    .A(_0393_));
 sg13g2_xnor2_1 _1238_ (.Y(_0499_),
    .A(_0393_),
    .B(_0497_));
 sg13g2_nor2_2 _1239_ (.A(_0396_),
    .B(_0412_),
    .Y(_0500_));
 sg13g2_inv_1 _1240_ (.Y(_0501_),
    .A(_0500_));
 sg13g2_xnor2_1 _1241_ (.Y(_0502_),
    .A(_0396_),
    .B(_0412_));
 sg13g2_nand3_1 _1242_ (.B(_0006_),
    .C(_0361_),
    .A(net100),
    .Y(_0503_));
 sg13g2_xor2_1 _1243_ (.B(_0503_),
    .A(net109),
    .X(_0504_));
 sg13g2_nor2_1 _1244_ (.A(_0502_),
    .B(_0504_),
    .Y(_0505_));
 sg13g2_xor2_1 _1245_ (.B(_0504_),
    .A(_0502_),
    .X(_0506_));
 sg13g2_nand2_1 _1246_ (.Y(_0507_),
    .A(_0469_),
    .B(_0506_));
 sg13g2_xnor2_1 _1247_ (.Y(_0508_),
    .A(_0469_),
    .B(_0506_));
 sg13g2_xnor2_1 _1248_ (.Y(_0509_),
    .A(_0499_),
    .B(_0508_));
 sg13g2_nand2b_1 _1249_ (.Y(_0510_),
    .B(_0495_),
    .A_N(_0509_));
 sg13g2_xor2_1 _1250_ (.B(_0509_),
    .A(_0495_),
    .X(_0511_));
 sg13g2_xor2_1 _1251_ (.B(_0511_),
    .A(_0494_),
    .X(_0512_));
 sg13g2_nand2_1 _1252_ (.Y(_0513_),
    .A(_0491_),
    .B(_0512_));
 sg13g2_xnor2_1 _1253_ (.Y(_0514_),
    .A(_0491_),
    .B(_0512_));
 sg13g2_xor2_1 _1254_ (.B(_0514_),
    .A(_0455_),
    .X(_0515_));
 sg13g2_nor2b_1 _1255_ (.A(_0482_),
    .B_N(_0515_),
    .Y(_0516_));
 sg13g2_xnor2_1 _1256_ (.Y(_0517_),
    .A(_0482_),
    .B(_0515_));
 sg13g2_nand2_1 _1257_ (.Y(_0518_),
    .A(_0487_),
    .B(_0517_));
 sg13g2_xnor2_1 _1258_ (.Y(_0519_),
    .A(_0487_),
    .B(_0517_));
 sg13g2_a21oi_1 _1259_ (.A1(_0452_),
    .A2(_0488_),
    .Y(_0520_),
    .B1(_0485_));
 sg13g2_or2_1 _1260_ (.X(_0521_),
    .B(_0520_),
    .A(_0519_));
 sg13g2_nand2_1 _1261_ (.Y(_0522_),
    .A(net126),
    .B(_0521_));
 sg13g2_a21oi_1 _1262_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0028_),
    .B1(_0522_));
 sg13g2_o21ai_1 _1263_ (.B1(_0513_),
    .Y(_0523_),
    .A1(_0455_),
    .A2(_0514_));
 sg13g2_o21ai_1 _1264_ (.B1(_0510_),
    .Y(_0524_),
    .A1(_0494_),
    .A2(_0511_));
 sg13g2_a21o_1 _1265_ (.A2(_0498_),
    .A1(_0496_),
    .B1(_0373_),
    .X(_0525_));
 sg13g2_nand3_1 _1266_ (.B(_0496_),
    .C(_0498_),
    .A(_0373_),
    .Y(_0526_));
 sg13g2_nand2_1 _1267_ (.Y(_0527_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_o21ai_1 _1268_ (.B1(_0507_),
    .Y(_0528_),
    .A1(_0499_),
    .A2(_0508_));
 sg13g2_xnor2_1 _1269_ (.Y(_0529_),
    .A(_0429_),
    .B(_0500_));
 sg13g2_nor2_1 _1270_ (.A(_0408_),
    .B(_0529_),
    .Y(_0530_));
 sg13g2_xnor2_1 _1271_ (.Y(_0531_),
    .A(_0408_),
    .B(_0529_));
 sg13g2_nor2_2 _1272_ (.A(_0412_),
    .B(_0431_),
    .Y(_0532_));
 sg13g2_xor2_1 _1273_ (.B(_0431_),
    .A(_0412_),
    .X(_0533_));
 sg13g2_nand2_1 _1274_ (.Y(_0534_),
    .A(_0687_),
    .B(_0533_));
 sg13g2_xnor2_1 _1275_ (.Y(_0535_),
    .A(_0004_),
    .B(_0533_));
 sg13g2_nand2_1 _1276_ (.Y(_0536_),
    .A(_0505_),
    .B(_0535_));
 sg13g2_xnor2_1 _1277_ (.Y(_0537_),
    .A(_0505_),
    .B(_0535_));
 sg13g2_xor2_1 _1278_ (.B(_0537_),
    .A(_0531_),
    .X(_0538_));
 sg13g2_nand2_1 _1279_ (.Y(_0539_),
    .A(_0528_),
    .B(_0538_));
 sg13g2_xnor2_1 _1280_ (.Y(_0540_),
    .A(_0528_),
    .B(_0538_));
 sg13g2_xor2_1 _1281_ (.B(_0540_),
    .A(_0527_),
    .X(_0541_));
 sg13g2_nand2_1 _1282_ (.Y(_0542_),
    .A(_0524_),
    .B(_0541_));
 sg13g2_xnor2_1 _1283_ (.Y(_0543_),
    .A(_0524_),
    .B(_0541_));
 sg13g2_xor2_1 _1284_ (.B(_0543_),
    .A(_0492_),
    .X(_0544_));
 sg13g2_nand2_1 _1285_ (.Y(_0545_),
    .A(_0523_),
    .B(_0544_));
 sg13g2_xor2_1 _1286_ (.B(_0544_),
    .A(_0523_),
    .X(_0546_));
 sg13g2_or2_1 _1287_ (.X(_0547_),
    .B(_0546_),
    .A(_0516_));
 sg13g2_xnor2_1 _1288_ (.Y(_0548_),
    .A(_0516_),
    .B(_0546_));
 sg13g2_and3_1 _1289_ (.X(_0549_),
    .A(_0518_),
    .B(_0521_),
    .C(_0548_));
 sg13g2_a21oi_1 _1290_ (.A1(_0518_),
    .A2(_0521_),
    .Y(_0550_),
    .B1(_0548_));
 sg13g2_nor3_1 _1291_ (.A(_0690_),
    .B(_0549_),
    .C(_0550_),
    .Y(_0029_));
 sg13g2_o21ai_1 _1292_ (.B1(_0542_),
    .Y(_0551_),
    .A1(_0492_),
    .A2(_0543_));
 sg13g2_o21ai_1 _1293_ (.B1(_0539_),
    .Y(_0552_),
    .A1(_0527_),
    .A2(_0540_));
 sg13g2_a21oi_1 _1294_ (.A1(_0429_),
    .A2(_0500_),
    .Y(_0553_),
    .B1(_0530_));
 sg13g2_xnor2_1 _1295_ (.Y(_0554_),
    .A(net95),
    .B(_0380_));
 sg13g2_or2_1 _1296_ (.X(_0555_),
    .B(_0554_),
    .A(_0553_));
 sg13g2_xnor2_1 _1297_ (.Y(_0556_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_o21ai_1 _1298_ (.B1(_0536_),
    .Y(_0557_),
    .A1(_0531_),
    .A2(_0537_));
 sg13g2_nor2b_1 _1299_ (.A(_0464_),
    .B_N(_0532_),
    .Y(_0558_));
 sg13g2_xnor2_1 _1300_ (.Y(_0559_),
    .A(_0464_),
    .B(_0532_));
 sg13g2_xnor2_1 _1301_ (.Y(_0560_),
    .A(_0427_),
    .B(_0559_));
 sg13g2_nor2_1 _1302_ (.A(_0431_),
    .B(_0468_),
    .Y(_0561_));
 sg13g2_xnor2_1 _1303_ (.Y(_0562_),
    .A(_0431_),
    .B(_0467_));
 sg13g2_nand2_1 _1304_ (.Y(_0563_),
    .A(net107),
    .B(_0562_));
 sg13g2_xnor2_1 _1305_ (.Y(_0564_),
    .A(net107),
    .B(_0562_));
 sg13g2_or2_1 _1306_ (.X(_0565_),
    .B(_0564_),
    .A(_0534_));
 sg13g2_xnor2_1 _1307_ (.Y(_0566_),
    .A(_0534_),
    .B(_0564_));
 sg13g2_xnor2_1 _1308_ (.Y(_0567_),
    .A(_0560_),
    .B(_0566_));
 sg13g2_nand2b_1 _1309_ (.Y(_0568_),
    .B(_0557_),
    .A_N(_0567_));
 sg13g2_xor2_1 _1310_ (.B(_0567_),
    .A(_0557_),
    .X(_0569_));
 sg13g2_xor2_1 _1311_ (.B(_0569_),
    .A(_0556_),
    .X(_0570_));
 sg13g2_nand2_1 _1312_ (.Y(_0571_),
    .A(_0552_),
    .B(_0570_));
 sg13g2_xnor2_1 _1313_ (.Y(_0572_),
    .A(_0552_),
    .B(_0570_));
 sg13g2_xnor2_1 _1314_ (.Y(_0573_),
    .A(_0525_),
    .B(_0572_));
 sg13g2_nand2b_1 _1315_ (.Y(_0574_),
    .B(_0551_),
    .A_N(_0573_));
 sg13g2_xor2_1 _1316_ (.B(_0573_),
    .A(_0551_),
    .X(_0575_));
 sg13g2_nor2_1 _1317_ (.A(_0545_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_inv_1 _1318_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_xnor2_1 _1319_ (.Y(_0578_),
    .A(_0545_),
    .B(_0575_));
 sg13g2_a22oi_1 _1320_ (.Y(_0579_),
    .B1(_0546_),
    .B2(_0516_),
    .A2(_0517_),
    .A1(_0487_));
 sg13g2_o21ai_1 _1321_ (.B1(_0579_),
    .Y(_0580_),
    .A1(_0519_),
    .A2(_0520_));
 sg13g2_nand2_1 _1322_ (.Y(_0581_),
    .A(_0547_),
    .B(_0580_));
 sg13g2_o21ai_1 _1323_ (.B1(net126),
    .Y(_0582_),
    .A1(_0578_),
    .A2(_0581_));
 sg13g2_a21oi_1 _1324_ (.A1(_0578_),
    .A2(_0581_),
    .Y(_0030_),
    .B1(_0582_));
 sg13g2_o21ai_1 _1325_ (.B1(_0571_),
    .Y(_0583_),
    .A1(_0525_),
    .A2(_0572_));
 sg13g2_o21ai_1 _1326_ (.B1(_0568_),
    .Y(_0584_),
    .A1(_0556_),
    .A2(_0569_));
 sg13g2_a21oi_1 _1327_ (.A1(_0427_),
    .A2(_0559_),
    .Y(_0585_),
    .B1(_0558_));
 sg13g2_nand2b_1 _1328_ (.Y(_0586_),
    .B(_0389_),
    .A_N(_0585_));
 sg13g2_xor2_1 _1329_ (.B(_0585_),
    .A(_0389_),
    .X(_0587_));
 sg13g2_xnor2_1 _1330_ (.Y(_0588_),
    .A(_0382_),
    .B(_0587_));
 sg13g2_o21ai_1 _1331_ (.B1(_0565_),
    .Y(_0589_),
    .A1(_0560_),
    .A2(_0566_));
 sg13g2_nor2_1 _1332_ (.A(_0468_),
    .B(_0504_),
    .Y(_0590_));
 sg13g2_xnor2_1 _1333_ (.Y(_0591_),
    .A(_0467_),
    .B(_0504_));
 sg13g2_nand2_1 _1334_ (.Y(_0592_),
    .A(net105),
    .B(_0591_));
 sg13g2_xnor2_1 _1335_ (.Y(_0593_),
    .A(net105),
    .B(_0591_));
 sg13g2_or2_1 _1336_ (.X(_0594_),
    .B(_0593_),
    .A(_0563_));
 sg13g2_xor2_1 _1337_ (.B(_0593_),
    .A(_0563_),
    .X(_0595_));
 sg13g2_nor2b_1 _1338_ (.A(_0502_),
    .B_N(_0561_),
    .Y(_0596_));
 sg13g2_xnor2_1 _1339_ (.Y(_0597_),
    .A(_0502_),
    .B(_0561_));
 sg13g2_xnor2_1 _1340_ (.Y(_0598_),
    .A(_0462_),
    .B(_0597_));
 sg13g2_nand2_1 _1341_ (.Y(_0599_),
    .A(_0595_),
    .B(_0598_));
 sg13g2_xnor2_1 _1342_ (.Y(_0600_),
    .A(_0595_),
    .B(_0598_));
 sg13g2_nor2b_1 _1343_ (.A(_0600_),
    .B_N(_0589_),
    .Y(_0601_));
 sg13g2_xor2_1 _1344_ (.B(_0600_),
    .A(_0589_),
    .X(_0602_));
 sg13g2_nor2_1 _1345_ (.A(_0588_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xor2_1 _1346_ (.B(_0602_),
    .A(_0588_),
    .X(_0604_));
 sg13g2_nand2_1 _1347_ (.Y(_0605_),
    .A(_0584_),
    .B(_0604_));
 sg13g2_xnor2_1 _1348_ (.Y(_0606_),
    .A(_0584_),
    .B(_0604_));
 sg13g2_xor2_1 _1349_ (.B(_0606_),
    .A(_0555_),
    .X(_0607_));
 sg13g2_nand2_1 _1350_ (.Y(_0608_),
    .A(_0583_),
    .B(_0607_));
 sg13g2_xnor2_1 _1351_ (.Y(_0609_),
    .A(_0583_),
    .B(_0607_));
 sg13g2_nor2_1 _1352_ (.A(_0574_),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_nand2_1 _1353_ (.Y(_0611_),
    .A(_0574_),
    .B(_0609_));
 sg13g2_xor2_1 _1354_ (.B(_0609_),
    .A(_0574_),
    .X(_0612_));
 sg13g2_o21ai_1 _1355_ (.B1(_0577_),
    .Y(_0613_),
    .A1(_0578_),
    .A2(_0581_));
 sg13g2_o21ai_1 _1356_ (.B1(net126),
    .Y(_0614_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_a21oi_1 _1357_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0031_),
    .B1(_0614_));
 sg13g2_nand2b_1 _1358_ (.Y(_0615_),
    .B(_0612_),
    .A_N(_0578_));
 sg13g2_nand3b_1 _1359_ (.B(_0580_),
    .C(_0547_),
    .Y(_0616_),
    .A_N(_0615_));
 sg13g2_a21oi_1 _1360_ (.A1(_0576_),
    .A2(_0611_),
    .Y(_0617_),
    .B1(_0610_));
 sg13g2_o21ai_1 _1361_ (.B1(_0586_),
    .Y(_0618_),
    .A1(_0382_),
    .A2(_0587_));
 sg13g2_nand2_1 _1362_ (.Y(_0619_),
    .A(_0358_),
    .B(_0618_));
 sg13g2_xor2_1 _1363_ (.B(_0618_),
    .A(_0358_),
    .X(_0620_));
 sg13g2_nor2_1 _1364_ (.A(_0601_),
    .B(_0603_),
    .Y(_0621_));
 sg13g2_nor2_1 _1365_ (.A(_0004_),
    .B(_0504_),
    .Y(_0622_));
 sg13g2_xnor2_1 _1366_ (.Y(_0623_),
    .A(_0687_),
    .B(_0504_));
 sg13g2_nand2_1 _1367_ (.Y(_0624_),
    .A(net100),
    .B(_0623_));
 sg13g2_xnor2_1 _1368_ (.Y(_0625_),
    .A(net100),
    .B(_0623_));
 sg13g2_xor2_1 _1369_ (.B(_0625_),
    .A(_0592_),
    .X(_0626_));
 sg13g2_nand2_1 _1370_ (.Y(_0627_),
    .A(_0533_),
    .B(_0590_));
 sg13g2_xnor2_1 _1371_ (.Y(_0628_),
    .A(_0533_),
    .B(_0590_));
 sg13g2_xnor2_1 _1372_ (.Y(_0629_),
    .A(_0500_),
    .B(_0628_));
 sg13g2_nand2_1 _1373_ (.Y(_0630_),
    .A(_0626_),
    .B(_0629_));
 sg13g2_xnor2_1 _1374_ (.Y(_0631_),
    .A(_0626_),
    .B(_0629_));
 sg13g2_a21oi_1 _1375_ (.A1(_0594_),
    .A2(_0599_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_nand3_1 _1376_ (.B(_0599_),
    .C(_0631_),
    .A(_0594_),
    .Y(_0633_));
 sg13g2_nand2b_1 _1377_ (.Y(_0634_),
    .B(_0633_),
    .A_N(_0632_));
 sg13g2_a21o_1 _1378_ (.A2(_0597_),
    .A1(_0461_),
    .B1(_0596_),
    .X(_0635_));
 sg13g2_xnor2_1 _1379_ (.Y(_0636_),
    .A(net95),
    .B(_0374_));
 sg13g2_nor2_1 _1380_ (.A(_0368_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_xor2_1 _1381_ (.B(_0636_),
    .A(_0368_),
    .X(_0638_));
 sg13g2_nand2_1 _1382_ (.Y(_0639_),
    .A(_0635_),
    .B(_0638_));
 sg13g2_xnor2_1 _1383_ (.Y(_0640_),
    .A(_0635_),
    .B(_0638_));
 sg13g2_xor2_1 _1384_ (.B(_0640_),
    .A(_0388_),
    .X(_0641_));
 sg13g2_nor2b_1 _1385_ (.A(_0634_),
    .B_N(_0641_),
    .Y(_0642_));
 sg13g2_xnor2_1 _1386_ (.Y(_0643_),
    .A(_0634_),
    .B(_0641_));
 sg13g2_nor2b_1 _1387_ (.A(_0621_),
    .B_N(_0643_),
    .Y(_0644_));
 sg13g2_xnor2_1 _1388_ (.Y(_0645_),
    .A(_0621_),
    .B(_0643_));
 sg13g2_xnor2_1 _1389_ (.Y(_0646_),
    .A(_0620_),
    .B(_0645_));
 sg13g2_o21ai_1 _1390_ (.B1(_0605_),
    .Y(_0647_),
    .A1(_0555_),
    .A2(_0606_));
 sg13g2_nor2b_1 _1391_ (.A(_0646_),
    .B_N(_0647_),
    .Y(_0648_));
 sg13g2_xor2_1 _1392_ (.B(_0647_),
    .A(_0646_),
    .X(_0649_));
 sg13g2_or2_1 _1393_ (.X(_0650_),
    .B(_0649_),
    .A(_0608_));
 sg13g2_xnor2_1 _1394_ (.Y(_0651_),
    .A(_0608_),
    .B(_0649_));
 sg13g2_nand3_1 _1395_ (.B(_0617_),
    .C(_0651_),
    .A(_0616_),
    .Y(_0652_));
 sg13g2_a21o_1 _1396_ (.A2(_0617_),
    .A1(_0616_),
    .B1(_0651_),
    .X(_0653_));
 sg13g2_and3_1 _1397_ (.X(_0032_),
    .A(net126),
    .B(_0652_),
    .C(_0653_));
 sg13g2_a21oi_1 _1398_ (.A1(_0620_),
    .A2(_0645_),
    .Y(_0654_),
    .B1(_0644_));
 sg13g2_o21ai_1 _1399_ (.B1(_0627_),
    .Y(_0655_),
    .A1(_0501_),
    .A2(_0628_));
 sg13g2_xnor2_1 _1400_ (.Y(_0656_),
    .A(_0399_),
    .B(_0655_));
 sg13g2_xnor2_1 _1401_ (.Y(_0657_),
    .A(_0689_),
    .B(_0237_));
 sg13g2_xnor2_1 _1402_ (.Y(_0658_),
    .A(_0357_),
    .B(_0657_));
 sg13g2_xnor2_1 _1403_ (.Y(_0659_),
    .A(_0562_),
    .B(_0622_));
 sg13g2_xnor2_1 _1404_ (.Y(_0660_),
    .A(_0532_),
    .B(_0624_));
 sg13g2_xnor2_1 _1405_ (.Y(_0661_),
    .A(_0658_),
    .B(_0660_));
 sg13g2_xnor2_1 _1406_ (.Y(_0662_),
    .A(_0659_),
    .B(_0661_));
 sg13g2_xnor2_1 _1407_ (.Y(_0663_),
    .A(_0656_),
    .B(_0662_));
 sg13g2_o21ai_1 _1408_ (.B1(_0630_),
    .Y(_0664_),
    .A1(_0592_),
    .A2(_0625_));
 sg13g2_xor2_1 _1409_ (.B(_0664_),
    .A(_0637_),
    .X(_0665_));
 sg13g2_xor2_1 _1410_ (.B(_0665_),
    .A(_0663_),
    .X(_0666_));
 sg13g2_o21ai_1 _1411_ (.B1(_0401_),
    .Y(_0667_),
    .A1(net95),
    .A2(_0374_));
 sg13g2_nor2_1 _1412_ (.A(_0632_),
    .B(_0642_),
    .Y(_0668_));
 sg13g2_o21ai_1 _1413_ (.B1(_0639_),
    .Y(_0669_),
    .A1(_0388_),
    .A2(_0640_));
 sg13g2_xor2_1 _1414_ (.B(_0669_),
    .A(_0667_),
    .X(_0670_));
 sg13g2_xnor2_1 _1415_ (.Y(_0671_),
    .A(_0666_),
    .B(_0670_));
 sg13g2_xnor2_1 _1416_ (.Y(_0672_),
    .A(_0668_),
    .B(_0671_));
 sg13g2_xnor2_1 _1417_ (.Y(_0673_),
    .A(_0654_),
    .B(_0672_));
 sg13g2_xnor2_1 _1418_ (.Y(_0674_),
    .A(_0619_),
    .B(_0648_));
 sg13g2_xnor2_1 _1419_ (.Y(_0675_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_a21oi_1 _1420_ (.A1(_0650_),
    .A2(_0653_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_and3_1 _1421_ (.X(_0677_),
    .A(_0650_),
    .B(_0653_),
    .C(_0675_));
 sg13g2_nor3_1 _1422_ (.A(_0690_),
    .B(_0676_),
    .C(_0677_),
    .Y(_0033_));
 sg13g2_dfrbp_1 _1423_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net32),
    .D(_0010_),
    .Q_N(_0009_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _1424_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net31),
    .D(_0011_),
    .Q_N(_0002_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1425_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net30),
    .D(_0012_),
    .Q_N(_0008_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1426_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net53),
    .D(_0013_),
    .Q_N(_0706_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _1427_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net52),
    .D(_0014_),
    .Q_N(_0007_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _1428_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net51),
    .D(_0015_),
    .Q_N(_0705_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 _1429_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net50),
    .D(_0016_),
    .Q_N(_0000_),
    .Q(\state[6] ));
 sg13g2_dfrbp_1 _1430_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net49),
    .D(_0017_),
    .Q_N(_0704_),
    .Q(\state[7] ));
 sg13g2_dfrbp_1 _1431_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(_0018_),
    .Q_N(_0001_),
    .Q(\state[8] ));
 sg13g2_dfrbp_1 _1432_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net47),
    .D(_0019_),
    .Q_N(_0003_),
    .Q(\state[9] ));
 sg13g2_dfrbp_1 _1433_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net46),
    .D(_0020_),
    .Q_N(_0703_),
    .Q(\state[10] ));
 sg13g2_dfrbp_1 _1434_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net45),
    .D(_0021_),
    .Q_N(_0004_),
    .Q(\state[11] ));
 sg13g2_dfrbp_1 _1435_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net44),
    .D(_0022_),
    .Q_N(_0702_),
    .Q(\state[12] ));
 sg13g2_dfrbp_1 _1436_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net43),
    .D(_0023_),
    .Q_N(_0701_),
    .Q(\state[13] ));
 sg13g2_dfrbp_1 _1437_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net42),
    .D(_0024_),
    .Q_N(_0005_),
    .Q(\state[14] ));
 sg13g2_dfrbp_1 _1438_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net41),
    .D(_0025_),
    .Q_N(_0006_),
    .Q(\state[15] ));
 sg13g2_dfrbp_1 _1439_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net40),
    .D(_0026_),
    .Q_N(_0700_),
    .Q(\pcg_out[0] ));
 sg13g2_dfrbp_1 _1440_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net39),
    .D(_0027_),
    .Q_N(_0699_),
    .Q(\pcg_out[1] ));
 sg13g2_dfrbp_1 _1441_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net38),
    .D(_0028_),
    .Q_N(_0698_),
    .Q(\pcg_out[2] ));
 sg13g2_dfrbp_1 _1442_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net37),
    .D(_0029_),
    .Q_N(_0697_),
    .Q(\pcg_out[3] ));
 sg13g2_dfrbp_1 _1443_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(_0030_),
    .Q_N(_0696_),
    .Q(\pcg_out[4] ));
 sg13g2_dfrbp_1 _1444_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(_0031_),
    .Q_N(_0695_),
    .Q(\pcg_out[5] ));
 sg13g2_dfrbp_1 _1445_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net34),
    .D(_0032_),
    .Q_N(_0694_),
    .Q(\pcg_out[6] ));
 sg13g2_dfrbp_1 _1446_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0033_),
    .Q_N(_0693_),
    .Q(\pcg_out[7] ));
 sg13g2_tiehi _1424__31 (.L_HI(net31));
 sg13g2_tiehi _1423__32 (.L_HI(net32));
 sg13g2_tiehi _1446__33 (.L_HI(net33));
 sg13g2_tiehi _1445__34 (.L_HI(net34));
 sg13g2_tiehi _1444__35 (.L_HI(net35));
 sg13g2_tiehi _1443__36 (.L_HI(net36));
 sg13g2_tiehi _1442__37 (.L_HI(net37));
 sg13g2_tiehi _1441__38 (.L_HI(net38));
 sg13g2_tiehi _1440__39 (.L_HI(net39));
 sg13g2_tiehi _1439__40 (.L_HI(net40));
 sg13g2_tiehi _1438__41 (.L_HI(net41));
 sg13g2_tiehi _1437__42 (.L_HI(net42));
 sg13g2_tiehi _1436__43 (.L_HI(net43));
 sg13g2_tiehi _1435__44 (.L_HI(net44));
 sg13g2_tiehi _1434__45 (.L_HI(net45));
 sg13g2_tiehi _1433__46 (.L_HI(net46));
 sg13g2_tiehi _1432__47 (.L_HI(net47));
 sg13g2_tiehi _1431__48 (.L_HI(net48));
 sg13g2_tiehi _1430__49 (.L_HI(net49));
 sg13g2_tiehi _1429__50 (.L_HI(net50));
 sg13g2_tiehi _1428__51 (.L_HI(net51));
 sg13g2_tiehi _1427__52 (.L_HI(net52));
 sg13g2_tiehi _1426__53 (.L_HI(net53));
 sg13g2_tiehi tt_um_crispy_vga_54 (.L_HI(net54));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_crispy_vga_17 (.L_LO(net17));
 sg13g2_tielo tt_um_crispy_vga_18 (.L_LO(net18));
 sg13g2_tielo tt_um_crispy_vga_19 (.L_LO(net19));
 sg13g2_tielo tt_um_crispy_vga_20 (.L_LO(net20));
 sg13g2_tielo tt_um_crispy_vga_21 (.L_LO(net21));
 sg13g2_tielo tt_um_crispy_vga_22 (.L_LO(net22));
 sg13g2_tielo tt_um_crispy_vga_23 (.L_LO(net23));
 sg13g2_tielo tt_um_crispy_vga_24 (.L_LO(net24));
 sg13g2_tielo tt_um_crispy_vga_25 (.L_LO(net25));
 sg13g2_tielo tt_um_crispy_vga_26 (.L_LO(net26));
 sg13g2_tielo tt_um_crispy_vga_27 (.L_LO(net27));
 sg13g2_tielo tt_um_crispy_vga_28 (.L_LO(net28));
 sg13g2_tielo tt_um_crispy_vga_29 (.L_LO(net29));
 sg13g2_tiehi _1425__30 (.L_HI(net30));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(_0350_));
 sg13g2_buf_2 fanout96 (.A(\state[15] ),
    .X(net96));
 sg13g2_buf_4 fanout97 (.X(net97),
    .A(net99));
 sg13g2_buf_1 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net100),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(\state[14] ),
    .X(net100));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net102));
 sg13g2_buf_1 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(\state[13] ),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(\state[12] ),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(\state[12] ),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(\state[11] ),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(\state[10] ),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(\state[10] ),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(\state[9] ),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(\state[8] ),
    .X(net112));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(\state[7] ));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(\state[6] ));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net116));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(\state[5] ));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(\state[4] ));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(\state[3] ));
 sg13g2_buf_1 fanout119 (.A(\state[3] ),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(\state[2] ));
 sg13g2_buf_2 fanout121 (.A(\state[1] ),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(\state[0] ),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net126));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(rst_n),
    .X(net126));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_tielo tt_um_crispy_vga_16 (.L_LO(net16));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0009_),
    .X(net55));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_decap_8 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_decap_8 FILLER_9_187 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_decap_8 FILLER_9_236 ();
 sg13g2_decap_8 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_250 ();
 sg13g2_decap_8 FILLER_9_257 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_285 ();
 sg13g2_decap_8 FILLER_9_292 ();
 sg13g2_decap_8 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_306 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_decap_4 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_decap_4 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_decap_4 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_decap_4 FILLER_11_107 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_127 ();
 sg13g2_fill_2 FILLER_11_134 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_157 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_4 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_2 FILLER_12_85 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_fill_2 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_178 ();
 sg13g2_fill_2 FILLER_12_206 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_decap_4 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_4 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_250 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_decap_8 FILLER_12_264 ();
 sg13g2_decap_8 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_278 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_114 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_152 ();
 sg13g2_decap_4 FILLER_13_159 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_decap_8 FILLER_13_170 ();
 sg13g2_fill_2 FILLER_13_177 ();
 sg13g2_decap_4 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_211 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_4 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_decap_4 FILLER_14_68 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_1 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_decap_4 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_176 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_93 ();
 sg13g2_fill_2 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_decap_4 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_159 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_fill_2 FILLER_15_211 ();
 sg13g2_decap_4 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_230 ();
 sg13g2_decap_4 FILLER_15_237 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_decap_4 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_94 ();
 sg13g2_decap_4 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_decap_4 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_decap_4 FILLER_17_139 ();
 sg13g2_decap_4 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_4 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_225 ();
 sg13g2_decap_4 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_decap_4 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_decap_4 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_54 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_4 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_162 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_240 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_decap_4 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_decap_4 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_4 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_33 ();
 sg13g2_fill_1 FILLER_19_40 ();
 sg13g2_fill_1 FILLER_19_65 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_decap_4 FILLER_19_129 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_decap_4 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_4 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_311 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_decap_8 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_decap_4 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_4 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_149 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_4 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_342 ();
 sg13g2_decap_4 FILLER_20_348 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_decap_4 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_fill_2 FILLER_21_80 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_decap_4 FILLER_21_96 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_4 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_decap_4 FILLER_22_337 ();
 sg13g2_decap_4 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_23 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_125 ();
 sg13g2_decap_4 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_fill_2 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_decap_4 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_decap_4 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_2 FILLER_24_59 ();
 sg13g2_fill_1 FILLER_24_61 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_61 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_72 ();
 sg13g2_decap_4 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_decap_4 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_decap_4 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_decap_4 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_decap_4 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_61 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_4 FILLER_26_214 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_115 ();
 sg13g2_decap_4 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_decap_4 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_decap_4 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_4 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_decap_8 FILLER_28_64 ();
 sg13g2_fill_2 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_73 ();
 sg13g2_decap_8 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_decap_4 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_decap_4 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_47 ();
 sg13g2_decap_4 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_142 ();
 sg13g2_decap_4 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_decap_4 FILLER_29_378 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_decap_8 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_decap_4 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_decap_8 FILLER_30_303 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_4 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_fill_2 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_138 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_266 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_354 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_4 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_4 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_325 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_decap_4 FILLER_36_389 ();
 sg13g2_fill_2 FILLER_36_393 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net16;
 assign uio_oe[1] = net17;
 assign uio_oe[2] = net18;
 assign uio_oe[3] = net19;
 assign uio_oe[4] = net20;
 assign uio_oe[5] = net21;
 assign uio_oe[6] = net22;
 assign uio_oe[7] = net54;
 assign uio_out[0] = net23;
 assign uio_out[1] = net24;
 assign uio_out[2] = net25;
 assign uio_out[3] = net26;
 assign uio_out[4] = net27;
 assign uio_out[5] = net28;
 assign uio_out[6] = net29;
endmodule

module tt_um_algofoogle_tt09_ring_osc3 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire dummy;
 wire osc;
 wire \tapped_ring.b0 ;
 wire \tapped_ring.b1 ;
 wire \tapped_ring.b1001 ;
 wire \tapped_ring.b101 ;
 wire \tapped_ring.b11 ;
 wire \tapped_ring.b21 ;
 wire \tapped_ring.b301 ;
 wire \tapped_ring.b31 ;
 wire \tapped_ring.b41 ;
 wire \tapped_ring.b51 ;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire \tapped_ring.c0/ins[1] ;
 wire \tapped_ring.c0/ins[2] ;
 wire \tapped_ring.c0/ins[3] ;
 wire \tapped_ring.c0/ins[4] ;
 wire \tapped_ring.c0/ins[5] ;
 wire \tapped_ring.c0/ins[6] ;
 wire \tapped_ring.c0/ins[7] ;
 wire \tapped_ring.c0/ins[8] ;
 wire \tapped_ring.c0/ins[9] ;
 wire \tapped_ring.c1/ins[1] ;
 wire \tapped_ring.c1/ins[2] ;
 wire \tapped_ring.c1/ins[3] ;
 wire \tapped_ring.c1/ins[4] ;
 wire \tapped_ring.c1/ins[5] ;
 wire \tapped_ring.c1/ins[6] ;
 wire \tapped_ring.c1/ins[7] ;
 wire \tapped_ring.c1/ins[8] ;
 wire \tapped_ring.c1/ins[9] ;
 wire \tapped_ring.c2/ins[1] ;
 wire \tapped_ring.c2/ins[2] ;
 wire \tapped_ring.c2/ins[3] ;
 wire \tapped_ring.c2/ins[4] ;
 wire \tapped_ring.c2/ins[5] ;
 wire \tapped_ring.c2/ins[6] ;
 wire \tapped_ring.c2/ins[7] ;
 wire \tapped_ring.c2/ins[8] ;
 wire \tapped_ring.c2/ins[9] ;
 wire \tapped_ring.c3/ins[1] ;
 wire \tapped_ring.c3/ins[2] ;
 wire \tapped_ring.c3/ins[3] ;
 wire \tapped_ring.c3/ins[4] ;
 wire \tapped_ring.c3/ins[5] ;
 wire \tapped_ring.c3/ins[6] ;
 wire \tapped_ring.c3/ins[7] ;
 wire \tapped_ring.c3/ins[8] ;
 wire \tapped_ring.c3/ins[9] ;
 wire \tapped_ring.c4/ins[1] ;
 wire \tapped_ring.c4/ins[2] ;
 wire \tapped_ring.c4/ins[3] ;
 wire \tapped_ring.c4/ins[4] ;
 wire \tapped_ring.c4/ins[5] ;
 wire \tapped_ring.c4/ins[6] ;
 wire \tapped_ring.c4/ins[7] ;
 wire \tapped_ring.c4/ins[8] ;
 wire \tapped_ring.c4/ins[9] ;
 wire \tapped_ring.c5/ins[10] ;
 wire \tapped_ring.c5/ins[11] ;
 wire \tapped_ring.c5/ins[12] ;
 wire \tapped_ring.c5/ins[13] ;
 wire \tapped_ring.c5/ins[14] ;
 wire \tapped_ring.c5/ins[15] ;
 wire \tapped_ring.c5/ins[16] ;
 wire \tapped_ring.c5/ins[17] ;
 wire \tapped_ring.c5/ins[18] ;
 wire \tapped_ring.c5/ins[19] ;
 wire \tapped_ring.c5/ins[1] ;
 wire \tapped_ring.c5/ins[20] ;
 wire \tapped_ring.c5/ins[21] ;
 wire \tapped_ring.c5/ins[22] ;
 wire \tapped_ring.c5/ins[23] ;
 wire \tapped_ring.c5/ins[24] ;
 wire \tapped_ring.c5/ins[25] ;
 wire \tapped_ring.c5/ins[26] ;
 wire \tapped_ring.c5/ins[27] ;
 wire \tapped_ring.c5/ins[28] ;
 wire \tapped_ring.c5/ins[29] ;
 wire \tapped_ring.c5/ins[2] ;
 wire \tapped_ring.c5/ins[30] ;
 wire \tapped_ring.c5/ins[31] ;
 wire \tapped_ring.c5/ins[32] ;
 wire \tapped_ring.c5/ins[33] ;
 wire \tapped_ring.c5/ins[34] ;
 wire \tapped_ring.c5/ins[35] ;
 wire \tapped_ring.c5/ins[36] ;
 wire \tapped_ring.c5/ins[37] ;
 wire \tapped_ring.c5/ins[38] ;
 wire \tapped_ring.c5/ins[39] ;
 wire \tapped_ring.c5/ins[3] ;
 wire \tapped_ring.c5/ins[40] ;
 wire \tapped_ring.c5/ins[41] ;
 wire \tapped_ring.c5/ins[42] ;
 wire \tapped_ring.c5/ins[43] ;
 wire \tapped_ring.c5/ins[44] ;
 wire \tapped_ring.c5/ins[45] ;
 wire \tapped_ring.c5/ins[46] ;
 wire \tapped_ring.c5/ins[47] ;
 wire \tapped_ring.c5/ins[48] ;
 wire \tapped_ring.c5/ins[49] ;
 wire \tapped_ring.c5/ins[4] ;
 wire \tapped_ring.c5/ins[5] ;
 wire \tapped_ring.c5/ins[6] ;
 wire \tapped_ring.c5/ins[7] ;
 wire \tapped_ring.c5/ins[8] ;
 wire \tapped_ring.c5/ins[9] ;
 wire \tapped_ring.c6/ins[100] ;
 wire \tapped_ring.c6/ins[101] ;
 wire \tapped_ring.c6/ins[102] ;
 wire \tapped_ring.c6/ins[103] ;
 wire \tapped_ring.c6/ins[104] ;
 wire \tapped_ring.c6/ins[105] ;
 wire \tapped_ring.c6/ins[106] ;
 wire \tapped_ring.c6/ins[107] ;
 wire \tapped_ring.c6/ins[108] ;
 wire \tapped_ring.c6/ins[109] ;
 wire \tapped_ring.c6/ins[10] ;
 wire \tapped_ring.c6/ins[110] ;
 wire \tapped_ring.c6/ins[111] ;
 wire \tapped_ring.c6/ins[112] ;
 wire \tapped_ring.c6/ins[113] ;
 wire \tapped_ring.c6/ins[114] ;
 wire \tapped_ring.c6/ins[115] ;
 wire \tapped_ring.c6/ins[116] ;
 wire \tapped_ring.c6/ins[117] ;
 wire \tapped_ring.c6/ins[118] ;
 wire \tapped_ring.c6/ins[119] ;
 wire \tapped_ring.c6/ins[11] ;
 wire \tapped_ring.c6/ins[120] ;
 wire \tapped_ring.c6/ins[121] ;
 wire \tapped_ring.c6/ins[122] ;
 wire \tapped_ring.c6/ins[123] ;
 wire \tapped_ring.c6/ins[124] ;
 wire \tapped_ring.c6/ins[125] ;
 wire \tapped_ring.c6/ins[126] ;
 wire \tapped_ring.c6/ins[127] ;
 wire \tapped_ring.c6/ins[128] ;
 wire \tapped_ring.c6/ins[129] ;
 wire \tapped_ring.c6/ins[12] ;
 wire \tapped_ring.c6/ins[130] ;
 wire \tapped_ring.c6/ins[131] ;
 wire \tapped_ring.c6/ins[132] ;
 wire \tapped_ring.c6/ins[133] ;
 wire \tapped_ring.c6/ins[134] ;
 wire \tapped_ring.c6/ins[135] ;
 wire \tapped_ring.c6/ins[136] ;
 wire \tapped_ring.c6/ins[137] ;
 wire \tapped_ring.c6/ins[138] ;
 wire \tapped_ring.c6/ins[139] ;
 wire \tapped_ring.c6/ins[13] ;
 wire \tapped_ring.c6/ins[140] ;
 wire \tapped_ring.c6/ins[141] ;
 wire \tapped_ring.c6/ins[142] ;
 wire \tapped_ring.c6/ins[143] ;
 wire \tapped_ring.c6/ins[144] ;
 wire \tapped_ring.c6/ins[145] ;
 wire \tapped_ring.c6/ins[146] ;
 wire \tapped_ring.c6/ins[147] ;
 wire \tapped_ring.c6/ins[148] ;
 wire \tapped_ring.c6/ins[149] ;
 wire \tapped_ring.c6/ins[14] ;
 wire \tapped_ring.c6/ins[150] ;
 wire \tapped_ring.c6/ins[151] ;
 wire \tapped_ring.c6/ins[152] ;
 wire \tapped_ring.c6/ins[153] ;
 wire \tapped_ring.c6/ins[154] ;
 wire \tapped_ring.c6/ins[155] ;
 wire \tapped_ring.c6/ins[156] ;
 wire \tapped_ring.c6/ins[157] ;
 wire \tapped_ring.c6/ins[158] ;
 wire \tapped_ring.c6/ins[159] ;
 wire \tapped_ring.c6/ins[15] ;
 wire \tapped_ring.c6/ins[160] ;
 wire \tapped_ring.c6/ins[161] ;
 wire \tapped_ring.c6/ins[162] ;
 wire \tapped_ring.c6/ins[163] ;
 wire \tapped_ring.c6/ins[164] ;
 wire \tapped_ring.c6/ins[165] ;
 wire \tapped_ring.c6/ins[166] ;
 wire \tapped_ring.c6/ins[167] ;
 wire \tapped_ring.c6/ins[168] ;
 wire \tapped_ring.c6/ins[169] ;
 wire \tapped_ring.c6/ins[16] ;
 wire \tapped_ring.c6/ins[170] ;
 wire \tapped_ring.c6/ins[171] ;
 wire \tapped_ring.c6/ins[172] ;
 wire \tapped_ring.c6/ins[173] ;
 wire \tapped_ring.c6/ins[174] ;
 wire \tapped_ring.c6/ins[175] ;
 wire \tapped_ring.c6/ins[176] ;
 wire \tapped_ring.c6/ins[177] ;
 wire \tapped_ring.c6/ins[178] ;
 wire \tapped_ring.c6/ins[179] ;
 wire \tapped_ring.c6/ins[17] ;
 wire \tapped_ring.c6/ins[180] ;
 wire \tapped_ring.c6/ins[181] ;
 wire \tapped_ring.c6/ins[182] ;
 wire \tapped_ring.c6/ins[183] ;
 wire \tapped_ring.c6/ins[184] ;
 wire \tapped_ring.c6/ins[185] ;
 wire \tapped_ring.c6/ins[186] ;
 wire \tapped_ring.c6/ins[187] ;
 wire \tapped_ring.c6/ins[188] ;
 wire \tapped_ring.c6/ins[189] ;
 wire \tapped_ring.c6/ins[18] ;
 wire \tapped_ring.c6/ins[190] ;
 wire \tapped_ring.c6/ins[191] ;
 wire \tapped_ring.c6/ins[192] ;
 wire \tapped_ring.c6/ins[193] ;
 wire \tapped_ring.c6/ins[194] ;
 wire \tapped_ring.c6/ins[195] ;
 wire \tapped_ring.c6/ins[196] ;
 wire \tapped_ring.c6/ins[197] ;
 wire \tapped_ring.c6/ins[198] ;
 wire \tapped_ring.c6/ins[199] ;
 wire \tapped_ring.c6/ins[19] ;
 wire \tapped_ring.c6/ins[1] ;
 wire \tapped_ring.c6/ins[20] ;
 wire \tapped_ring.c6/ins[21] ;
 wire \tapped_ring.c6/ins[22] ;
 wire \tapped_ring.c6/ins[23] ;
 wire \tapped_ring.c6/ins[24] ;
 wire \tapped_ring.c6/ins[25] ;
 wire \tapped_ring.c6/ins[26] ;
 wire \tapped_ring.c6/ins[27] ;
 wire \tapped_ring.c6/ins[28] ;
 wire \tapped_ring.c6/ins[29] ;
 wire \tapped_ring.c6/ins[2] ;
 wire \tapped_ring.c6/ins[30] ;
 wire \tapped_ring.c6/ins[31] ;
 wire \tapped_ring.c6/ins[32] ;
 wire \tapped_ring.c6/ins[33] ;
 wire \tapped_ring.c6/ins[34] ;
 wire \tapped_ring.c6/ins[35] ;
 wire \tapped_ring.c6/ins[36] ;
 wire \tapped_ring.c6/ins[37] ;
 wire \tapped_ring.c6/ins[38] ;
 wire \tapped_ring.c6/ins[39] ;
 wire \tapped_ring.c6/ins[3] ;
 wire \tapped_ring.c6/ins[40] ;
 wire \tapped_ring.c6/ins[41] ;
 wire \tapped_ring.c6/ins[42] ;
 wire \tapped_ring.c6/ins[43] ;
 wire \tapped_ring.c6/ins[44] ;
 wire \tapped_ring.c6/ins[45] ;
 wire \tapped_ring.c6/ins[46] ;
 wire \tapped_ring.c6/ins[47] ;
 wire \tapped_ring.c6/ins[48] ;
 wire \tapped_ring.c6/ins[49] ;
 wire \tapped_ring.c6/ins[4] ;
 wire \tapped_ring.c6/ins[50] ;
 wire \tapped_ring.c6/ins[51] ;
 wire \tapped_ring.c6/ins[52] ;
 wire \tapped_ring.c6/ins[53] ;
 wire \tapped_ring.c6/ins[54] ;
 wire \tapped_ring.c6/ins[55] ;
 wire \tapped_ring.c6/ins[56] ;
 wire \tapped_ring.c6/ins[57] ;
 wire \tapped_ring.c6/ins[58] ;
 wire \tapped_ring.c6/ins[59] ;
 wire \tapped_ring.c6/ins[5] ;
 wire \tapped_ring.c6/ins[60] ;
 wire \tapped_ring.c6/ins[61] ;
 wire \tapped_ring.c6/ins[62] ;
 wire \tapped_ring.c6/ins[63] ;
 wire \tapped_ring.c6/ins[64] ;
 wire \tapped_ring.c6/ins[65] ;
 wire \tapped_ring.c6/ins[66] ;
 wire \tapped_ring.c6/ins[67] ;
 wire \tapped_ring.c6/ins[68] ;
 wire \tapped_ring.c6/ins[69] ;
 wire \tapped_ring.c6/ins[6] ;
 wire \tapped_ring.c6/ins[70] ;
 wire \tapped_ring.c6/ins[71] ;
 wire \tapped_ring.c6/ins[72] ;
 wire \tapped_ring.c6/ins[73] ;
 wire \tapped_ring.c6/ins[74] ;
 wire \tapped_ring.c6/ins[75] ;
 wire \tapped_ring.c6/ins[76] ;
 wire \tapped_ring.c6/ins[77] ;
 wire \tapped_ring.c6/ins[78] ;
 wire \tapped_ring.c6/ins[79] ;
 wire \tapped_ring.c6/ins[7] ;
 wire \tapped_ring.c6/ins[80] ;
 wire \tapped_ring.c6/ins[81] ;
 wire \tapped_ring.c6/ins[82] ;
 wire \tapped_ring.c6/ins[83] ;
 wire \tapped_ring.c6/ins[84] ;
 wire \tapped_ring.c6/ins[85] ;
 wire \tapped_ring.c6/ins[86] ;
 wire \tapped_ring.c6/ins[87] ;
 wire \tapped_ring.c6/ins[88] ;
 wire \tapped_ring.c6/ins[89] ;
 wire \tapped_ring.c6/ins[8] ;
 wire \tapped_ring.c6/ins[90] ;
 wire \tapped_ring.c6/ins[91] ;
 wire \tapped_ring.c6/ins[92] ;
 wire \tapped_ring.c6/ins[93] ;
 wire \tapped_ring.c6/ins[94] ;
 wire \tapped_ring.c6/ins[95] ;
 wire \tapped_ring.c6/ins[96] ;
 wire \tapped_ring.c6/ins[97] ;
 wire \tapped_ring.c6/ins[98] ;
 wire \tapped_ring.c6/ins[99] ;
 wire \tapped_ring.c6/ins[9] ;
 wire \tapped_ring.c7/ins[100] ;
 wire \tapped_ring.c7/ins[101] ;
 wire \tapped_ring.c7/ins[102] ;
 wire \tapped_ring.c7/ins[103] ;
 wire \tapped_ring.c7/ins[104] ;
 wire \tapped_ring.c7/ins[105] ;
 wire \tapped_ring.c7/ins[106] ;
 wire \tapped_ring.c7/ins[107] ;
 wire \tapped_ring.c7/ins[108] ;
 wire \tapped_ring.c7/ins[109] ;
 wire \tapped_ring.c7/ins[10] ;
 wire \tapped_ring.c7/ins[110] ;
 wire \tapped_ring.c7/ins[111] ;
 wire \tapped_ring.c7/ins[112] ;
 wire \tapped_ring.c7/ins[113] ;
 wire \tapped_ring.c7/ins[114] ;
 wire \tapped_ring.c7/ins[115] ;
 wire \tapped_ring.c7/ins[116] ;
 wire \tapped_ring.c7/ins[117] ;
 wire \tapped_ring.c7/ins[118] ;
 wire \tapped_ring.c7/ins[119] ;
 wire \tapped_ring.c7/ins[11] ;
 wire \tapped_ring.c7/ins[120] ;
 wire \tapped_ring.c7/ins[121] ;
 wire \tapped_ring.c7/ins[122] ;
 wire \tapped_ring.c7/ins[123] ;
 wire \tapped_ring.c7/ins[124] ;
 wire \tapped_ring.c7/ins[125] ;
 wire \tapped_ring.c7/ins[126] ;
 wire \tapped_ring.c7/ins[127] ;
 wire \tapped_ring.c7/ins[128] ;
 wire \tapped_ring.c7/ins[129] ;
 wire \tapped_ring.c7/ins[12] ;
 wire \tapped_ring.c7/ins[130] ;
 wire \tapped_ring.c7/ins[131] ;
 wire \tapped_ring.c7/ins[132] ;
 wire \tapped_ring.c7/ins[133] ;
 wire \tapped_ring.c7/ins[134] ;
 wire \tapped_ring.c7/ins[135] ;
 wire \tapped_ring.c7/ins[136] ;
 wire \tapped_ring.c7/ins[137] ;
 wire \tapped_ring.c7/ins[138] ;
 wire \tapped_ring.c7/ins[139] ;
 wire \tapped_ring.c7/ins[13] ;
 wire \tapped_ring.c7/ins[140] ;
 wire \tapped_ring.c7/ins[141] ;
 wire \tapped_ring.c7/ins[142] ;
 wire \tapped_ring.c7/ins[143] ;
 wire \tapped_ring.c7/ins[144] ;
 wire \tapped_ring.c7/ins[145] ;
 wire \tapped_ring.c7/ins[146] ;
 wire \tapped_ring.c7/ins[147] ;
 wire \tapped_ring.c7/ins[148] ;
 wire \tapped_ring.c7/ins[149] ;
 wire \tapped_ring.c7/ins[14] ;
 wire \tapped_ring.c7/ins[150] ;
 wire \tapped_ring.c7/ins[151] ;
 wire \tapped_ring.c7/ins[152] ;
 wire \tapped_ring.c7/ins[153] ;
 wire \tapped_ring.c7/ins[154] ;
 wire \tapped_ring.c7/ins[155] ;
 wire \tapped_ring.c7/ins[156] ;
 wire \tapped_ring.c7/ins[157] ;
 wire \tapped_ring.c7/ins[158] ;
 wire \tapped_ring.c7/ins[159] ;
 wire \tapped_ring.c7/ins[15] ;
 wire \tapped_ring.c7/ins[160] ;
 wire \tapped_ring.c7/ins[161] ;
 wire \tapped_ring.c7/ins[162] ;
 wire \tapped_ring.c7/ins[163] ;
 wire \tapped_ring.c7/ins[164] ;
 wire \tapped_ring.c7/ins[165] ;
 wire \tapped_ring.c7/ins[166] ;
 wire \tapped_ring.c7/ins[167] ;
 wire \tapped_ring.c7/ins[168] ;
 wire \tapped_ring.c7/ins[169] ;
 wire \tapped_ring.c7/ins[16] ;
 wire \tapped_ring.c7/ins[170] ;
 wire \tapped_ring.c7/ins[171] ;
 wire \tapped_ring.c7/ins[172] ;
 wire \tapped_ring.c7/ins[173] ;
 wire \tapped_ring.c7/ins[174] ;
 wire \tapped_ring.c7/ins[175] ;
 wire \tapped_ring.c7/ins[176] ;
 wire \tapped_ring.c7/ins[177] ;
 wire \tapped_ring.c7/ins[178] ;
 wire \tapped_ring.c7/ins[179] ;
 wire \tapped_ring.c7/ins[17] ;
 wire \tapped_ring.c7/ins[180] ;
 wire \tapped_ring.c7/ins[181] ;
 wire \tapped_ring.c7/ins[182] ;
 wire \tapped_ring.c7/ins[183] ;
 wire \tapped_ring.c7/ins[184] ;
 wire \tapped_ring.c7/ins[185] ;
 wire \tapped_ring.c7/ins[186] ;
 wire \tapped_ring.c7/ins[187] ;
 wire \tapped_ring.c7/ins[188] ;
 wire \tapped_ring.c7/ins[189] ;
 wire \tapped_ring.c7/ins[18] ;
 wire \tapped_ring.c7/ins[190] ;
 wire \tapped_ring.c7/ins[191] ;
 wire \tapped_ring.c7/ins[192] ;
 wire \tapped_ring.c7/ins[193] ;
 wire \tapped_ring.c7/ins[194] ;
 wire \tapped_ring.c7/ins[195] ;
 wire \tapped_ring.c7/ins[196] ;
 wire \tapped_ring.c7/ins[197] ;
 wire \tapped_ring.c7/ins[198] ;
 wire \tapped_ring.c7/ins[199] ;
 wire \tapped_ring.c7/ins[19] ;
 wire \tapped_ring.c7/ins[1] ;
 wire \tapped_ring.c7/ins[200] ;
 wire \tapped_ring.c7/ins[201] ;
 wire \tapped_ring.c7/ins[202] ;
 wire \tapped_ring.c7/ins[203] ;
 wire \tapped_ring.c7/ins[204] ;
 wire \tapped_ring.c7/ins[205] ;
 wire \tapped_ring.c7/ins[206] ;
 wire \tapped_ring.c7/ins[207] ;
 wire \tapped_ring.c7/ins[208] ;
 wire \tapped_ring.c7/ins[209] ;
 wire \tapped_ring.c7/ins[20] ;
 wire \tapped_ring.c7/ins[210] ;
 wire \tapped_ring.c7/ins[211] ;
 wire \tapped_ring.c7/ins[212] ;
 wire \tapped_ring.c7/ins[213] ;
 wire \tapped_ring.c7/ins[214] ;
 wire \tapped_ring.c7/ins[215] ;
 wire \tapped_ring.c7/ins[216] ;
 wire \tapped_ring.c7/ins[217] ;
 wire \tapped_ring.c7/ins[218] ;
 wire \tapped_ring.c7/ins[219] ;
 wire \tapped_ring.c7/ins[21] ;
 wire \tapped_ring.c7/ins[220] ;
 wire \tapped_ring.c7/ins[221] ;
 wire \tapped_ring.c7/ins[222] ;
 wire \tapped_ring.c7/ins[223] ;
 wire \tapped_ring.c7/ins[224] ;
 wire \tapped_ring.c7/ins[225] ;
 wire \tapped_ring.c7/ins[226] ;
 wire \tapped_ring.c7/ins[227] ;
 wire \tapped_ring.c7/ins[228] ;
 wire \tapped_ring.c7/ins[229] ;
 wire \tapped_ring.c7/ins[22] ;
 wire \tapped_ring.c7/ins[230] ;
 wire \tapped_ring.c7/ins[231] ;
 wire \tapped_ring.c7/ins[232] ;
 wire \tapped_ring.c7/ins[233] ;
 wire \tapped_ring.c7/ins[234] ;
 wire \tapped_ring.c7/ins[235] ;
 wire \tapped_ring.c7/ins[236] ;
 wire \tapped_ring.c7/ins[237] ;
 wire \tapped_ring.c7/ins[238] ;
 wire \tapped_ring.c7/ins[239] ;
 wire \tapped_ring.c7/ins[23] ;
 wire \tapped_ring.c7/ins[240] ;
 wire \tapped_ring.c7/ins[241] ;
 wire \tapped_ring.c7/ins[242] ;
 wire \tapped_ring.c7/ins[243] ;
 wire \tapped_ring.c7/ins[244] ;
 wire \tapped_ring.c7/ins[245] ;
 wire \tapped_ring.c7/ins[246] ;
 wire \tapped_ring.c7/ins[247] ;
 wire \tapped_ring.c7/ins[248] ;
 wire \tapped_ring.c7/ins[249] ;
 wire \tapped_ring.c7/ins[24] ;
 wire \tapped_ring.c7/ins[250] ;
 wire \tapped_ring.c7/ins[251] ;
 wire \tapped_ring.c7/ins[252] ;
 wire \tapped_ring.c7/ins[253] ;
 wire \tapped_ring.c7/ins[254] ;
 wire \tapped_ring.c7/ins[255] ;
 wire \tapped_ring.c7/ins[256] ;
 wire \tapped_ring.c7/ins[257] ;
 wire \tapped_ring.c7/ins[258] ;
 wire \tapped_ring.c7/ins[259] ;
 wire \tapped_ring.c7/ins[25] ;
 wire \tapped_ring.c7/ins[260] ;
 wire \tapped_ring.c7/ins[261] ;
 wire \tapped_ring.c7/ins[262] ;
 wire \tapped_ring.c7/ins[263] ;
 wire \tapped_ring.c7/ins[264] ;
 wire \tapped_ring.c7/ins[265] ;
 wire \tapped_ring.c7/ins[266] ;
 wire \tapped_ring.c7/ins[267] ;
 wire \tapped_ring.c7/ins[268] ;
 wire \tapped_ring.c7/ins[269] ;
 wire \tapped_ring.c7/ins[26] ;
 wire \tapped_ring.c7/ins[270] ;
 wire \tapped_ring.c7/ins[271] ;
 wire \tapped_ring.c7/ins[272] ;
 wire \tapped_ring.c7/ins[273] ;
 wire \tapped_ring.c7/ins[274] ;
 wire \tapped_ring.c7/ins[275] ;
 wire \tapped_ring.c7/ins[276] ;
 wire \tapped_ring.c7/ins[277] ;
 wire \tapped_ring.c7/ins[278] ;
 wire \tapped_ring.c7/ins[279] ;
 wire \tapped_ring.c7/ins[27] ;
 wire \tapped_ring.c7/ins[280] ;
 wire \tapped_ring.c7/ins[281] ;
 wire \tapped_ring.c7/ins[282] ;
 wire \tapped_ring.c7/ins[283] ;
 wire \tapped_ring.c7/ins[284] ;
 wire \tapped_ring.c7/ins[285] ;
 wire \tapped_ring.c7/ins[286] ;
 wire \tapped_ring.c7/ins[287] ;
 wire \tapped_ring.c7/ins[288] ;
 wire \tapped_ring.c7/ins[289] ;
 wire \tapped_ring.c7/ins[28] ;
 wire \tapped_ring.c7/ins[290] ;
 wire \tapped_ring.c7/ins[291] ;
 wire \tapped_ring.c7/ins[292] ;
 wire \tapped_ring.c7/ins[293] ;
 wire \tapped_ring.c7/ins[294] ;
 wire \tapped_ring.c7/ins[295] ;
 wire \tapped_ring.c7/ins[296] ;
 wire \tapped_ring.c7/ins[297] ;
 wire \tapped_ring.c7/ins[298] ;
 wire \tapped_ring.c7/ins[299] ;
 wire \tapped_ring.c7/ins[29] ;
 wire \tapped_ring.c7/ins[2] ;
 wire \tapped_ring.c7/ins[300] ;
 wire \tapped_ring.c7/ins[301] ;
 wire \tapped_ring.c7/ins[302] ;
 wire \tapped_ring.c7/ins[303] ;
 wire \tapped_ring.c7/ins[304] ;
 wire \tapped_ring.c7/ins[305] ;
 wire \tapped_ring.c7/ins[306] ;
 wire \tapped_ring.c7/ins[307] ;
 wire \tapped_ring.c7/ins[308] ;
 wire \tapped_ring.c7/ins[309] ;
 wire \tapped_ring.c7/ins[30] ;
 wire \tapped_ring.c7/ins[310] ;
 wire \tapped_ring.c7/ins[311] ;
 wire \tapped_ring.c7/ins[312] ;
 wire \tapped_ring.c7/ins[313] ;
 wire \tapped_ring.c7/ins[314] ;
 wire \tapped_ring.c7/ins[315] ;
 wire \tapped_ring.c7/ins[316] ;
 wire \tapped_ring.c7/ins[317] ;
 wire \tapped_ring.c7/ins[318] ;
 wire \tapped_ring.c7/ins[319] ;
 wire \tapped_ring.c7/ins[31] ;
 wire \tapped_ring.c7/ins[320] ;
 wire \tapped_ring.c7/ins[321] ;
 wire \tapped_ring.c7/ins[322] ;
 wire \tapped_ring.c7/ins[323] ;
 wire \tapped_ring.c7/ins[324] ;
 wire \tapped_ring.c7/ins[325] ;
 wire \tapped_ring.c7/ins[326] ;
 wire \tapped_ring.c7/ins[327] ;
 wire \tapped_ring.c7/ins[328] ;
 wire \tapped_ring.c7/ins[329] ;
 wire \tapped_ring.c7/ins[32] ;
 wire \tapped_ring.c7/ins[330] ;
 wire \tapped_ring.c7/ins[331] ;
 wire \tapped_ring.c7/ins[332] ;
 wire \tapped_ring.c7/ins[333] ;
 wire \tapped_ring.c7/ins[334] ;
 wire \tapped_ring.c7/ins[335] ;
 wire \tapped_ring.c7/ins[336] ;
 wire \tapped_ring.c7/ins[337] ;
 wire \tapped_ring.c7/ins[338] ;
 wire \tapped_ring.c7/ins[339] ;
 wire \tapped_ring.c7/ins[33] ;
 wire \tapped_ring.c7/ins[340] ;
 wire \tapped_ring.c7/ins[341] ;
 wire \tapped_ring.c7/ins[342] ;
 wire \tapped_ring.c7/ins[343] ;
 wire \tapped_ring.c7/ins[344] ;
 wire \tapped_ring.c7/ins[345] ;
 wire \tapped_ring.c7/ins[346] ;
 wire \tapped_ring.c7/ins[347] ;
 wire \tapped_ring.c7/ins[348] ;
 wire \tapped_ring.c7/ins[349] ;
 wire \tapped_ring.c7/ins[34] ;
 wire \tapped_ring.c7/ins[350] ;
 wire \tapped_ring.c7/ins[351] ;
 wire \tapped_ring.c7/ins[352] ;
 wire \tapped_ring.c7/ins[353] ;
 wire \tapped_ring.c7/ins[354] ;
 wire \tapped_ring.c7/ins[355] ;
 wire \tapped_ring.c7/ins[356] ;
 wire \tapped_ring.c7/ins[357] ;
 wire \tapped_ring.c7/ins[358] ;
 wire \tapped_ring.c7/ins[359] ;
 wire \tapped_ring.c7/ins[35] ;
 wire \tapped_ring.c7/ins[360] ;
 wire \tapped_ring.c7/ins[361] ;
 wire \tapped_ring.c7/ins[362] ;
 wire \tapped_ring.c7/ins[363] ;
 wire \tapped_ring.c7/ins[364] ;
 wire \tapped_ring.c7/ins[365] ;
 wire \tapped_ring.c7/ins[366] ;
 wire \tapped_ring.c7/ins[367] ;
 wire \tapped_ring.c7/ins[368] ;
 wire \tapped_ring.c7/ins[369] ;
 wire \tapped_ring.c7/ins[36] ;
 wire \tapped_ring.c7/ins[370] ;
 wire \tapped_ring.c7/ins[371] ;
 wire \tapped_ring.c7/ins[372] ;
 wire \tapped_ring.c7/ins[373] ;
 wire \tapped_ring.c7/ins[374] ;
 wire \tapped_ring.c7/ins[375] ;
 wire \tapped_ring.c7/ins[376] ;
 wire \tapped_ring.c7/ins[377] ;
 wire \tapped_ring.c7/ins[378] ;
 wire \tapped_ring.c7/ins[379] ;
 wire \tapped_ring.c7/ins[37] ;
 wire \tapped_ring.c7/ins[380] ;
 wire \tapped_ring.c7/ins[381] ;
 wire \tapped_ring.c7/ins[382] ;
 wire \tapped_ring.c7/ins[383] ;
 wire \tapped_ring.c7/ins[384] ;
 wire \tapped_ring.c7/ins[385] ;
 wire \tapped_ring.c7/ins[386] ;
 wire \tapped_ring.c7/ins[387] ;
 wire \tapped_ring.c7/ins[388] ;
 wire \tapped_ring.c7/ins[389] ;
 wire \tapped_ring.c7/ins[38] ;
 wire \tapped_ring.c7/ins[390] ;
 wire \tapped_ring.c7/ins[391] ;
 wire \tapped_ring.c7/ins[392] ;
 wire \tapped_ring.c7/ins[393] ;
 wire \tapped_ring.c7/ins[394] ;
 wire \tapped_ring.c7/ins[395] ;
 wire \tapped_ring.c7/ins[396] ;
 wire \tapped_ring.c7/ins[397] ;
 wire \tapped_ring.c7/ins[398] ;
 wire \tapped_ring.c7/ins[399] ;
 wire \tapped_ring.c7/ins[39] ;
 wire \tapped_ring.c7/ins[3] ;
 wire \tapped_ring.c7/ins[400] ;
 wire \tapped_ring.c7/ins[401] ;
 wire \tapped_ring.c7/ins[402] ;
 wire \tapped_ring.c7/ins[403] ;
 wire \tapped_ring.c7/ins[404] ;
 wire \tapped_ring.c7/ins[405] ;
 wire \tapped_ring.c7/ins[406] ;
 wire \tapped_ring.c7/ins[407] ;
 wire \tapped_ring.c7/ins[408] ;
 wire \tapped_ring.c7/ins[409] ;
 wire \tapped_ring.c7/ins[40] ;
 wire \tapped_ring.c7/ins[410] ;
 wire \tapped_ring.c7/ins[411] ;
 wire \tapped_ring.c7/ins[412] ;
 wire \tapped_ring.c7/ins[413] ;
 wire \tapped_ring.c7/ins[414] ;
 wire \tapped_ring.c7/ins[415] ;
 wire \tapped_ring.c7/ins[416] ;
 wire \tapped_ring.c7/ins[417] ;
 wire \tapped_ring.c7/ins[418] ;
 wire \tapped_ring.c7/ins[419] ;
 wire \tapped_ring.c7/ins[41] ;
 wire \tapped_ring.c7/ins[420] ;
 wire \tapped_ring.c7/ins[421] ;
 wire \tapped_ring.c7/ins[422] ;
 wire \tapped_ring.c7/ins[423] ;
 wire \tapped_ring.c7/ins[424] ;
 wire \tapped_ring.c7/ins[425] ;
 wire \tapped_ring.c7/ins[426] ;
 wire \tapped_ring.c7/ins[427] ;
 wire \tapped_ring.c7/ins[428] ;
 wire \tapped_ring.c7/ins[429] ;
 wire \tapped_ring.c7/ins[42] ;
 wire \tapped_ring.c7/ins[430] ;
 wire \tapped_ring.c7/ins[431] ;
 wire \tapped_ring.c7/ins[432] ;
 wire \tapped_ring.c7/ins[433] ;
 wire \tapped_ring.c7/ins[434] ;
 wire \tapped_ring.c7/ins[435] ;
 wire \tapped_ring.c7/ins[436] ;
 wire \tapped_ring.c7/ins[437] ;
 wire \tapped_ring.c7/ins[438] ;
 wire \tapped_ring.c7/ins[439] ;
 wire \tapped_ring.c7/ins[43] ;
 wire \tapped_ring.c7/ins[440] ;
 wire \tapped_ring.c7/ins[441] ;
 wire \tapped_ring.c7/ins[442] ;
 wire \tapped_ring.c7/ins[443] ;
 wire \tapped_ring.c7/ins[444] ;
 wire \tapped_ring.c7/ins[445] ;
 wire \tapped_ring.c7/ins[446] ;
 wire \tapped_ring.c7/ins[447] ;
 wire \tapped_ring.c7/ins[448] ;
 wire \tapped_ring.c7/ins[449] ;
 wire \tapped_ring.c7/ins[44] ;
 wire \tapped_ring.c7/ins[450] ;
 wire \tapped_ring.c7/ins[451] ;
 wire \tapped_ring.c7/ins[452] ;
 wire \tapped_ring.c7/ins[453] ;
 wire \tapped_ring.c7/ins[454] ;
 wire \tapped_ring.c7/ins[455] ;
 wire \tapped_ring.c7/ins[456] ;
 wire \tapped_ring.c7/ins[457] ;
 wire \tapped_ring.c7/ins[458] ;
 wire \tapped_ring.c7/ins[459] ;
 wire \tapped_ring.c7/ins[45] ;
 wire \tapped_ring.c7/ins[460] ;
 wire \tapped_ring.c7/ins[461] ;
 wire \tapped_ring.c7/ins[462] ;
 wire \tapped_ring.c7/ins[463] ;
 wire \tapped_ring.c7/ins[464] ;
 wire \tapped_ring.c7/ins[465] ;
 wire \tapped_ring.c7/ins[466] ;
 wire \tapped_ring.c7/ins[467] ;
 wire \tapped_ring.c7/ins[468] ;
 wire \tapped_ring.c7/ins[469] ;
 wire \tapped_ring.c7/ins[46] ;
 wire \tapped_ring.c7/ins[470] ;
 wire \tapped_ring.c7/ins[471] ;
 wire \tapped_ring.c7/ins[472] ;
 wire \tapped_ring.c7/ins[473] ;
 wire \tapped_ring.c7/ins[474] ;
 wire \tapped_ring.c7/ins[475] ;
 wire \tapped_ring.c7/ins[476] ;
 wire \tapped_ring.c7/ins[477] ;
 wire \tapped_ring.c7/ins[478] ;
 wire \tapped_ring.c7/ins[479] ;
 wire \tapped_ring.c7/ins[47] ;
 wire \tapped_ring.c7/ins[480] ;
 wire \tapped_ring.c7/ins[481] ;
 wire \tapped_ring.c7/ins[482] ;
 wire \tapped_ring.c7/ins[483] ;
 wire \tapped_ring.c7/ins[484] ;
 wire \tapped_ring.c7/ins[485] ;
 wire \tapped_ring.c7/ins[486] ;
 wire \tapped_ring.c7/ins[487] ;
 wire \tapped_ring.c7/ins[488] ;
 wire \tapped_ring.c7/ins[489] ;
 wire \tapped_ring.c7/ins[48] ;
 wire \tapped_ring.c7/ins[490] ;
 wire \tapped_ring.c7/ins[491] ;
 wire \tapped_ring.c7/ins[492] ;
 wire \tapped_ring.c7/ins[493] ;
 wire \tapped_ring.c7/ins[494] ;
 wire \tapped_ring.c7/ins[495] ;
 wire \tapped_ring.c7/ins[496] ;
 wire \tapped_ring.c7/ins[497] ;
 wire \tapped_ring.c7/ins[498] ;
 wire \tapped_ring.c7/ins[499] ;
 wire \tapped_ring.c7/ins[49] ;
 wire \tapped_ring.c7/ins[4] ;
 wire \tapped_ring.c7/ins[500] ;
 wire \tapped_ring.c7/ins[501] ;
 wire \tapped_ring.c7/ins[502] ;
 wire \tapped_ring.c7/ins[503] ;
 wire \tapped_ring.c7/ins[504] ;
 wire \tapped_ring.c7/ins[505] ;
 wire \tapped_ring.c7/ins[506] ;
 wire \tapped_ring.c7/ins[507] ;
 wire \tapped_ring.c7/ins[508] ;
 wire \tapped_ring.c7/ins[509] ;
 wire \tapped_ring.c7/ins[50] ;
 wire \tapped_ring.c7/ins[510] ;
 wire \tapped_ring.c7/ins[511] ;
 wire \tapped_ring.c7/ins[512] ;
 wire \tapped_ring.c7/ins[513] ;
 wire \tapped_ring.c7/ins[514] ;
 wire \tapped_ring.c7/ins[515] ;
 wire \tapped_ring.c7/ins[516] ;
 wire \tapped_ring.c7/ins[517] ;
 wire \tapped_ring.c7/ins[518] ;
 wire \tapped_ring.c7/ins[519] ;
 wire \tapped_ring.c7/ins[51] ;
 wire \tapped_ring.c7/ins[520] ;
 wire \tapped_ring.c7/ins[521] ;
 wire \tapped_ring.c7/ins[522] ;
 wire \tapped_ring.c7/ins[523] ;
 wire \tapped_ring.c7/ins[524] ;
 wire \tapped_ring.c7/ins[525] ;
 wire \tapped_ring.c7/ins[526] ;
 wire \tapped_ring.c7/ins[527] ;
 wire \tapped_ring.c7/ins[528] ;
 wire \tapped_ring.c7/ins[529] ;
 wire \tapped_ring.c7/ins[52] ;
 wire \tapped_ring.c7/ins[530] ;
 wire \tapped_ring.c7/ins[531] ;
 wire \tapped_ring.c7/ins[532] ;
 wire \tapped_ring.c7/ins[533] ;
 wire \tapped_ring.c7/ins[534] ;
 wire \tapped_ring.c7/ins[535] ;
 wire \tapped_ring.c7/ins[536] ;
 wire \tapped_ring.c7/ins[537] ;
 wire \tapped_ring.c7/ins[538] ;
 wire \tapped_ring.c7/ins[539] ;
 wire \tapped_ring.c7/ins[53] ;
 wire \tapped_ring.c7/ins[540] ;
 wire \tapped_ring.c7/ins[541] ;
 wire \tapped_ring.c7/ins[542] ;
 wire \tapped_ring.c7/ins[543] ;
 wire \tapped_ring.c7/ins[544] ;
 wire \tapped_ring.c7/ins[545] ;
 wire \tapped_ring.c7/ins[546] ;
 wire \tapped_ring.c7/ins[547] ;
 wire \tapped_ring.c7/ins[548] ;
 wire \tapped_ring.c7/ins[549] ;
 wire \tapped_ring.c7/ins[54] ;
 wire \tapped_ring.c7/ins[550] ;
 wire \tapped_ring.c7/ins[551] ;
 wire \tapped_ring.c7/ins[552] ;
 wire \tapped_ring.c7/ins[553] ;
 wire \tapped_ring.c7/ins[554] ;
 wire \tapped_ring.c7/ins[555] ;
 wire \tapped_ring.c7/ins[556] ;
 wire \tapped_ring.c7/ins[557] ;
 wire \tapped_ring.c7/ins[558] ;
 wire \tapped_ring.c7/ins[559] ;
 wire \tapped_ring.c7/ins[55] ;
 wire \tapped_ring.c7/ins[560] ;
 wire \tapped_ring.c7/ins[561] ;
 wire \tapped_ring.c7/ins[562] ;
 wire \tapped_ring.c7/ins[563] ;
 wire \tapped_ring.c7/ins[564] ;
 wire \tapped_ring.c7/ins[565] ;
 wire \tapped_ring.c7/ins[566] ;
 wire \tapped_ring.c7/ins[567] ;
 wire \tapped_ring.c7/ins[568] ;
 wire \tapped_ring.c7/ins[569] ;
 wire \tapped_ring.c7/ins[56] ;
 wire \tapped_ring.c7/ins[570] ;
 wire \tapped_ring.c7/ins[571] ;
 wire \tapped_ring.c7/ins[572] ;
 wire \tapped_ring.c7/ins[573] ;
 wire \tapped_ring.c7/ins[574] ;
 wire \tapped_ring.c7/ins[575] ;
 wire \tapped_ring.c7/ins[576] ;
 wire \tapped_ring.c7/ins[577] ;
 wire \tapped_ring.c7/ins[578] ;
 wire \tapped_ring.c7/ins[579] ;
 wire \tapped_ring.c7/ins[57] ;
 wire \tapped_ring.c7/ins[580] ;
 wire \tapped_ring.c7/ins[581] ;
 wire \tapped_ring.c7/ins[582] ;
 wire \tapped_ring.c7/ins[583] ;
 wire \tapped_ring.c7/ins[584] ;
 wire \tapped_ring.c7/ins[585] ;
 wire \tapped_ring.c7/ins[586] ;
 wire \tapped_ring.c7/ins[587] ;
 wire \tapped_ring.c7/ins[588] ;
 wire \tapped_ring.c7/ins[589] ;
 wire \tapped_ring.c7/ins[58] ;
 wire \tapped_ring.c7/ins[590] ;
 wire \tapped_ring.c7/ins[591] ;
 wire \tapped_ring.c7/ins[592] ;
 wire \tapped_ring.c7/ins[593] ;
 wire \tapped_ring.c7/ins[594] ;
 wire \tapped_ring.c7/ins[595] ;
 wire \tapped_ring.c7/ins[596] ;
 wire \tapped_ring.c7/ins[597] ;
 wire \tapped_ring.c7/ins[598] ;
 wire \tapped_ring.c7/ins[599] ;
 wire \tapped_ring.c7/ins[59] ;
 wire \tapped_ring.c7/ins[5] ;
 wire \tapped_ring.c7/ins[600] ;
 wire \tapped_ring.c7/ins[601] ;
 wire \tapped_ring.c7/ins[602] ;
 wire \tapped_ring.c7/ins[603] ;
 wire \tapped_ring.c7/ins[604] ;
 wire \tapped_ring.c7/ins[605] ;
 wire \tapped_ring.c7/ins[606] ;
 wire \tapped_ring.c7/ins[607] ;
 wire \tapped_ring.c7/ins[608] ;
 wire \tapped_ring.c7/ins[609] ;
 wire \tapped_ring.c7/ins[60] ;
 wire \tapped_ring.c7/ins[610] ;
 wire \tapped_ring.c7/ins[611] ;
 wire \tapped_ring.c7/ins[612] ;
 wire \tapped_ring.c7/ins[613] ;
 wire \tapped_ring.c7/ins[614] ;
 wire \tapped_ring.c7/ins[615] ;
 wire \tapped_ring.c7/ins[616] ;
 wire \tapped_ring.c7/ins[617] ;
 wire \tapped_ring.c7/ins[618] ;
 wire \tapped_ring.c7/ins[619] ;
 wire \tapped_ring.c7/ins[61] ;
 wire \tapped_ring.c7/ins[620] ;
 wire \tapped_ring.c7/ins[621] ;
 wire \tapped_ring.c7/ins[622] ;
 wire \tapped_ring.c7/ins[623] ;
 wire \tapped_ring.c7/ins[624] ;
 wire \tapped_ring.c7/ins[625] ;
 wire \tapped_ring.c7/ins[626] ;
 wire \tapped_ring.c7/ins[627] ;
 wire \tapped_ring.c7/ins[628] ;
 wire \tapped_ring.c7/ins[629] ;
 wire \tapped_ring.c7/ins[62] ;
 wire \tapped_ring.c7/ins[630] ;
 wire \tapped_ring.c7/ins[631] ;
 wire \tapped_ring.c7/ins[632] ;
 wire \tapped_ring.c7/ins[633] ;
 wire \tapped_ring.c7/ins[634] ;
 wire \tapped_ring.c7/ins[635] ;
 wire \tapped_ring.c7/ins[636] ;
 wire \tapped_ring.c7/ins[637] ;
 wire \tapped_ring.c7/ins[638] ;
 wire \tapped_ring.c7/ins[639] ;
 wire \tapped_ring.c7/ins[63] ;
 wire \tapped_ring.c7/ins[640] ;
 wire \tapped_ring.c7/ins[641] ;
 wire \tapped_ring.c7/ins[642] ;
 wire \tapped_ring.c7/ins[643] ;
 wire \tapped_ring.c7/ins[644] ;
 wire \tapped_ring.c7/ins[645] ;
 wire \tapped_ring.c7/ins[646] ;
 wire \tapped_ring.c7/ins[647] ;
 wire \tapped_ring.c7/ins[648] ;
 wire \tapped_ring.c7/ins[649] ;
 wire \tapped_ring.c7/ins[64] ;
 wire \tapped_ring.c7/ins[650] ;
 wire \tapped_ring.c7/ins[651] ;
 wire \tapped_ring.c7/ins[652] ;
 wire \tapped_ring.c7/ins[653] ;
 wire \tapped_ring.c7/ins[654] ;
 wire \tapped_ring.c7/ins[655] ;
 wire \tapped_ring.c7/ins[656] ;
 wire \tapped_ring.c7/ins[657] ;
 wire \tapped_ring.c7/ins[658] ;
 wire \tapped_ring.c7/ins[659] ;
 wire \tapped_ring.c7/ins[65] ;
 wire \tapped_ring.c7/ins[660] ;
 wire \tapped_ring.c7/ins[661] ;
 wire \tapped_ring.c7/ins[662] ;
 wire \tapped_ring.c7/ins[663] ;
 wire \tapped_ring.c7/ins[664] ;
 wire \tapped_ring.c7/ins[665] ;
 wire \tapped_ring.c7/ins[666] ;
 wire \tapped_ring.c7/ins[667] ;
 wire \tapped_ring.c7/ins[668] ;
 wire \tapped_ring.c7/ins[669] ;
 wire \tapped_ring.c7/ins[66] ;
 wire \tapped_ring.c7/ins[670] ;
 wire \tapped_ring.c7/ins[671] ;
 wire \tapped_ring.c7/ins[672] ;
 wire \tapped_ring.c7/ins[673] ;
 wire \tapped_ring.c7/ins[674] ;
 wire \tapped_ring.c7/ins[675] ;
 wire \tapped_ring.c7/ins[676] ;
 wire \tapped_ring.c7/ins[677] ;
 wire \tapped_ring.c7/ins[678] ;
 wire \tapped_ring.c7/ins[679] ;
 wire \tapped_ring.c7/ins[67] ;
 wire \tapped_ring.c7/ins[680] ;
 wire \tapped_ring.c7/ins[681] ;
 wire \tapped_ring.c7/ins[682] ;
 wire \tapped_ring.c7/ins[683] ;
 wire \tapped_ring.c7/ins[684] ;
 wire \tapped_ring.c7/ins[685] ;
 wire \tapped_ring.c7/ins[686] ;
 wire \tapped_ring.c7/ins[687] ;
 wire \tapped_ring.c7/ins[688] ;
 wire \tapped_ring.c7/ins[689] ;
 wire \tapped_ring.c7/ins[68] ;
 wire \tapped_ring.c7/ins[690] ;
 wire \tapped_ring.c7/ins[691] ;
 wire \tapped_ring.c7/ins[692] ;
 wire \tapped_ring.c7/ins[693] ;
 wire \tapped_ring.c7/ins[694] ;
 wire \tapped_ring.c7/ins[695] ;
 wire \tapped_ring.c7/ins[696] ;
 wire \tapped_ring.c7/ins[697] ;
 wire \tapped_ring.c7/ins[698] ;
 wire \tapped_ring.c7/ins[699] ;
 wire \tapped_ring.c7/ins[69] ;
 wire \tapped_ring.c7/ins[6] ;
 wire \tapped_ring.c7/ins[70] ;
 wire \tapped_ring.c7/ins[71] ;
 wire \tapped_ring.c7/ins[72] ;
 wire \tapped_ring.c7/ins[73] ;
 wire \tapped_ring.c7/ins[74] ;
 wire \tapped_ring.c7/ins[75] ;
 wire \tapped_ring.c7/ins[76] ;
 wire \tapped_ring.c7/ins[77] ;
 wire \tapped_ring.c7/ins[78] ;
 wire \tapped_ring.c7/ins[79] ;
 wire \tapped_ring.c7/ins[7] ;
 wire \tapped_ring.c7/ins[80] ;
 wire \tapped_ring.c7/ins[81] ;
 wire \tapped_ring.c7/ins[82] ;
 wire \tapped_ring.c7/ins[83] ;
 wire \tapped_ring.c7/ins[84] ;
 wire \tapped_ring.c7/ins[85] ;
 wire \tapped_ring.c7/ins[86] ;
 wire \tapped_ring.c7/ins[87] ;
 wire \tapped_ring.c7/ins[88] ;
 wire \tapped_ring.c7/ins[89] ;
 wire \tapped_ring.c7/ins[8] ;
 wire \tapped_ring.c7/ins[90] ;
 wire \tapped_ring.c7/ins[91] ;
 wire \tapped_ring.c7/ins[92] ;
 wire \tapped_ring.c7/ins[93] ;
 wire \tapped_ring.c7/ins[94] ;
 wire \tapped_ring.c7/ins[95] ;
 wire \tapped_ring.c7/ins[96] ;
 wire \tapped_ring.c7/ins[97] ;
 wire \tapped_ring.c7/ins[98] ;
 wire \tapped_ring.c7/ins[99] ;
 wire \tapped_ring.c7/ins[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;

 sg13g2_inv_1 _38_ (.Y(_06_),
    .A(net4));
 sg13g2_inv_1 _39_ (.Y(_07_),
    .A(uo_out[4]));
 sg13g2_and4_1 _40_ (.A(net7),
    .B(net6),
    .C(net9),
    .D(net8),
    .X(_08_));
 sg13g2_nand3_1 _41_ (.B(net5),
    .C(_08_),
    .A(net4),
    .Y(_09_));
 sg13g2_nand4_1 _42_ (.B(net18),
    .C(net3),
    .A(net19),
    .Y(_10_),
    .D(net2));
 sg13g2_nand4_1 _43_ (.B(net14),
    .C(net17),
    .A(net15),
    .Y(_11_),
    .D(net16));
 sg13g2_nand4_1 _44_ (.B(net10),
    .C(net13),
    .A(net11),
    .Y(_12_),
    .D(net12));
 sg13g2_nor4_1 _45_ (.A(_09_),
    .B(_10_),
    .C(_11_),
    .D(_12_),
    .Y(dummy));
 sg13g2_mux2_1 _46_ (.A0(\tapped_ring.b31 ),
    .A1(\tapped_ring.b301 ),
    .S(net6),
    .X(_13_));
 sg13g2_nor2_1 _47_ (.A(net4),
    .B(_13_),
    .Y(_14_));
 sg13g2_mux2_1 _48_ (.A0(\tapped_ring.b41 ),
    .A1(\tapped_ring.b1001 ),
    .S(net6),
    .X(_15_));
 sg13g2_o21ai_1 _49_ (.B1(net5),
    .Y(_16_),
    .A1(_06_),
    .A2(_15_));
 sg13g2_mux4_1 _50_ (.S0(net4),
    .A0(\tapped_ring.b11 ),
    .A1(\tapped_ring.b21 ),
    .A2(\tapped_ring.b51 ),
    .A3(\tapped_ring.b101 ),
    .S1(net6),
    .X(_17_));
 sg13g2_nand2b_1 _51_ (.Y(_18_),
    .B(_17_),
    .A_N(net5));
 sg13g2_o21ai_1 _52_ (.B1(_18_),
    .Y(osc),
    .A1(_14_),
    .A2(_16_));
 sg13g2_and2_1 _53_ (.A(net2),
    .B(osc),
    .X(\tapped_ring.b0 ));
 sg13g2_xor2_1 _54_ (.B(uo_out[1]),
    .A(uo_out[2]),
    .X(_00_));
 sg13g2_nand3_1 _55_ (.B(uo_out[1]),
    .C(uo_out[3]),
    .A(uo_out[2]),
    .Y(_19_));
 sg13g2_a21o_1 _56_ (.A2(uo_out[1]),
    .A1(uo_out[2]),
    .B1(uo_out[3]),
    .X(_20_));
 sg13g2_and2_1 _57_ (.A(_19_),
    .B(_20_),
    .X(_01_));
 sg13g2_nor2_1 _58_ (.A(_07_),
    .B(_19_),
    .Y(_21_));
 sg13g2_xnor2_1 _59_ (.Y(_02_),
    .A(uo_out[4]),
    .B(_19_));
 sg13g2_xor2_1 _60_ (.B(_21_),
    .A(uo_out[5]),
    .X(_03_));
 sg13g2_nand3_1 _61_ (.B(uo_out[6]),
    .C(_21_),
    .A(uo_out[5]),
    .Y(_22_));
 sg13g2_a21o_1 _62_ (.A2(_21_),
    .A1(uo_out[5]),
    .B1(uo_out[6]),
    .X(_23_));
 sg13g2_and2_1 _63_ (.A(_22_),
    .B(_23_),
    .X(_04_));
 sg13g2_xnor2_1 _64_ (.Y(_05_),
    .A(uo_out[7]),
    .B(_22_));
 sg13g2_dfrbp_1 _65_ (.CLK(net1),
    .RESET_B(net36),
    .D(_24_),
    .Q_N(_24_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _66_ (.CLK(net1),
    .RESET_B(net37),
    .D(_00_),
    .Q_N(_26_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _67_ (.CLK(net1),
    .RESET_B(net38),
    .D(_01_),
    .Q_N(_27_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _68_ (.CLK(net1),
    .RESET_B(net39),
    .D(_02_),
    .Q_N(_28_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _69_ (.CLK(net1),
    .RESET_B(net40),
    .D(_03_),
    .Q_N(_29_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _70_ (.CLK(net1),
    .RESET_B(net34),
    .D(_04_),
    .Q_N(_30_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _71_ (.CLK(net1),
    .RESET_B(net35),
    .D(_05_),
    .Q_N(_25_),
    .Q(uo_out[7]));
 sg13g2_tiehi _71__34 (.L_HI(net35));
 sg13g2_tiehi _65__35 (.L_HI(net36));
 sg13g2_tiehi _66__36 (.L_HI(net37));
 sg13g2_tiehi _67__37 (.L_HI(net38));
 sg13g2_tiehi _68__38 (.L_HI(net39));
 sg13g2_tiehi _69__39 (.L_HI(net40));
 sg13g2_tiehi tt_um_algofoogle_tt09_ring_osc3_40 (.L_HI(net41));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_20 (.L_LO(net21));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_21 (.L_LO(net22));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_22 (.L_LO(net23));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_23 (.L_LO(net24));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_24 (.L_LO(net25));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_25 (.L_LO(net26));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_26 (.L_LO(net27));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_27 (.L_LO(net28));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_28 (.L_LO(net29));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_29 (.L_LO(net30));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_30 (.L_LO(net31));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_31 (.L_LO(net32));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_32 (.L_LO(net33));
 sg13g2_tiehi _70__33 (.L_HI(net34));
 sg13g2_buf_1 _94_ (.A(dummy),
    .X(uio_out[0]));
 sg13g2_buf_1 _95_ (.A(net1),
    .X(uo_out[0]));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[1] ),
    .A(\tapped_ring.b1 ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[2] ),
    .A(\tapped_ring.c0/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[3] ),
    .A(\tapped_ring.c0/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[4] ),
    .A(\tapped_ring.c0/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[5] ),
    .A(\tapped_ring.c0/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[6] ),
    .A(\tapped_ring.c0/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[7] ),
    .A(\tapped_ring.c0/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[8] ),
    .A(\tapped_ring.c0/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c0/ins[9] ),
    .A(\tapped_ring.c0/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c0/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.b11 ),
    .A(\tapped_ring.c0/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[1] ),
    .A(\tapped_ring.b11 ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[2] ),
    .A(\tapped_ring.c1/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[3] ),
    .A(\tapped_ring.c1/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[4] ),
    .A(\tapped_ring.c1/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[5] ),
    .A(\tapped_ring.c1/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[6] ),
    .A(\tapped_ring.c1/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[7] ),
    .A(\tapped_ring.c1/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[8] ),
    .A(\tapped_ring.c1/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c1/ins[9] ),
    .A(\tapped_ring.c1/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c1/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.b21 ),
    .A(\tapped_ring.c1/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[1] ),
    .A(\tapped_ring.b21 ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[2] ),
    .A(\tapped_ring.c2/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[3] ),
    .A(\tapped_ring.c2/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[4] ),
    .A(\tapped_ring.c2/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[5] ),
    .A(\tapped_ring.c2/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[6] ),
    .A(\tapped_ring.c2/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[7] ),
    .A(\tapped_ring.c2/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[8] ),
    .A(\tapped_ring.c2/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c2/ins[9] ),
    .A(\tapped_ring.c2/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c2/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.b31 ),
    .A(\tapped_ring.c2/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[1] ),
    .A(\tapped_ring.b31 ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[2] ),
    .A(\tapped_ring.c3/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[3] ),
    .A(\tapped_ring.c3/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[4] ),
    .A(\tapped_ring.c3/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[5] ),
    .A(\tapped_ring.c3/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[6] ),
    .A(\tapped_ring.c3/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[7] ),
    .A(\tapped_ring.c3/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[8] ),
    .A(\tapped_ring.c3/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c3/ins[9] ),
    .A(\tapped_ring.c3/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c3/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.b41 ),
    .A(\tapped_ring.c3/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[1] ),
    .A(\tapped_ring.b41 ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[2] ),
    .A(\tapped_ring.c4/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[3] ),
    .A(\tapped_ring.c4/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[4] ),
    .A(\tapped_ring.c4/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[5] ),
    .A(\tapped_ring.c4/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[6] ),
    .A(\tapped_ring.c4/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[7] ),
    .A(\tapped_ring.c4/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[8] ),
    .A(\tapped_ring.c4/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c4/ins[9] ),
    .A(\tapped_ring.c4/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c4/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.b51 ),
    .A(\tapped_ring.c4/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[1] ),
    .A(\tapped_ring.b51 ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[10]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[11] ),
    .A(\tapped_ring.c5/ins[10] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[11]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[12] ),
    .A(\tapped_ring.c5/ins[11] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[12]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[13] ),
    .A(\tapped_ring.c5/ins[12] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[13]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[14] ),
    .A(\tapped_ring.c5/ins[13] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[14]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[15] ),
    .A(\tapped_ring.c5/ins[14] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[15]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[16] ),
    .A(\tapped_ring.c5/ins[15] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[16]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[17] ),
    .A(\tapped_ring.c5/ins[16] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[17]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[18] ),
    .A(\tapped_ring.c5/ins[17] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[18]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[19] ),
    .A(\tapped_ring.c5/ins[18] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[19]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[20] ),
    .A(\tapped_ring.c5/ins[19] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[2] ),
    .A(\tapped_ring.c5/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[20]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[21] ),
    .A(\tapped_ring.c5/ins[20] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[21]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[22] ),
    .A(\tapped_ring.c5/ins[21] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[22]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[23] ),
    .A(\tapped_ring.c5/ins[22] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[23]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[24] ),
    .A(\tapped_ring.c5/ins[23] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[24]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[25] ),
    .A(\tapped_ring.c5/ins[24] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[25]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[26] ),
    .A(\tapped_ring.c5/ins[25] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[26]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[27] ),
    .A(\tapped_ring.c5/ins[26] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[27]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[28] ),
    .A(\tapped_ring.c5/ins[27] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[28]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[29] ),
    .A(\tapped_ring.c5/ins[28] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[29]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[30] ),
    .A(\tapped_ring.c5/ins[29] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[3] ),
    .A(\tapped_ring.c5/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[30]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[31] ),
    .A(\tapped_ring.c5/ins[30] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[31]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[32] ),
    .A(\tapped_ring.c5/ins[31] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[32]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[33] ),
    .A(\tapped_ring.c5/ins[32] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[33]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[34] ),
    .A(\tapped_ring.c5/ins[33] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[34]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[35] ),
    .A(\tapped_ring.c5/ins[34] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[35]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[36] ),
    .A(\tapped_ring.c5/ins[35] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[36]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[37] ),
    .A(\tapped_ring.c5/ins[36] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[37]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[38] ),
    .A(\tapped_ring.c5/ins[37] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[38]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[39] ),
    .A(\tapped_ring.c5/ins[38] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[39]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[40] ),
    .A(\tapped_ring.c5/ins[39] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[4] ),
    .A(\tapped_ring.c5/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[40]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[41] ),
    .A(\tapped_ring.c5/ins[40] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[41]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[42] ),
    .A(\tapped_ring.c5/ins[41] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[42]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[43] ),
    .A(\tapped_ring.c5/ins[42] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[43]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[44] ),
    .A(\tapped_ring.c5/ins[43] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[44]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[45] ),
    .A(\tapped_ring.c5/ins[44] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[45]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[46] ),
    .A(\tapped_ring.c5/ins[45] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[46]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[47] ),
    .A(\tapped_ring.c5/ins[46] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[47]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[48] ),
    .A(\tapped_ring.c5/ins[47] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[48]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[49] ),
    .A(\tapped_ring.c5/ins[48] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[49]/sky_inverter/_0_  (.Y(\tapped_ring.b101 ),
    .A(\tapped_ring.c5/ins[49] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[5] ),
    .A(\tapped_ring.c5/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[6] ),
    .A(\tapped_ring.c5/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[7] ),
    .A(\tapped_ring.c5/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[8] ),
    .A(\tapped_ring.c5/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[9] ),
    .A(\tapped_ring.c5/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c5/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.c5/ins[10] ),
    .A(\tapped_ring.c5/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[1] ),
    .A(\tapped_ring.b101 ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[100]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[101] ),
    .A(\tapped_ring.c6/ins[100] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[101]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[102] ),
    .A(\tapped_ring.c6/ins[101] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[102]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[103] ),
    .A(\tapped_ring.c6/ins[102] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[103]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[104] ),
    .A(\tapped_ring.c6/ins[103] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[104]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[105] ),
    .A(\tapped_ring.c6/ins[104] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[105]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[106] ),
    .A(\tapped_ring.c6/ins[105] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[106]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[107] ),
    .A(\tapped_ring.c6/ins[106] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[107]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[108] ),
    .A(\tapped_ring.c6/ins[107] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[108]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[109] ),
    .A(\tapped_ring.c6/ins[108] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[109]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[110] ),
    .A(\tapped_ring.c6/ins[109] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[10]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[11] ),
    .A(\tapped_ring.c6/ins[10] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[110]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[111] ),
    .A(\tapped_ring.c6/ins[110] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[111]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[112] ),
    .A(\tapped_ring.c6/ins[111] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[112]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[113] ),
    .A(\tapped_ring.c6/ins[112] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[113]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[114] ),
    .A(\tapped_ring.c6/ins[113] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[114]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[115] ),
    .A(\tapped_ring.c6/ins[114] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[115]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[116] ),
    .A(\tapped_ring.c6/ins[115] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[116]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[117] ),
    .A(\tapped_ring.c6/ins[116] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[117]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[118] ),
    .A(\tapped_ring.c6/ins[117] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[118]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[119] ),
    .A(\tapped_ring.c6/ins[118] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[119]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[120] ),
    .A(\tapped_ring.c6/ins[119] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[11]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[12] ),
    .A(\tapped_ring.c6/ins[11] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[120]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[121] ),
    .A(\tapped_ring.c6/ins[120] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[121]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[122] ),
    .A(\tapped_ring.c6/ins[121] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[122]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[123] ),
    .A(\tapped_ring.c6/ins[122] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[123]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[124] ),
    .A(\tapped_ring.c6/ins[123] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[124]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[125] ),
    .A(\tapped_ring.c6/ins[124] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[125]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[126] ),
    .A(\tapped_ring.c6/ins[125] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[126]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[127] ),
    .A(\tapped_ring.c6/ins[126] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[127]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[128] ),
    .A(\tapped_ring.c6/ins[127] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[128]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[129] ),
    .A(\tapped_ring.c6/ins[128] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[129]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[130] ),
    .A(\tapped_ring.c6/ins[129] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[12]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[13] ),
    .A(\tapped_ring.c6/ins[12] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[130]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[131] ),
    .A(\tapped_ring.c6/ins[130] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[131]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[132] ),
    .A(\tapped_ring.c6/ins[131] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[132]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[133] ),
    .A(\tapped_ring.c6/ins[132] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[133]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[134] ),
    .A(\tapped_ring.c6/ins[133] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[134]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[135] ),
    .A(\tapped_ring.c6/ins[134] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[135]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[136] ),
    .A(\tapped_ring.c6/ins[135] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[136]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[137] ),
    .A(\tapped_ring.c6/ins[136] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[137]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[138] ),
    .A(\tapped_ring.c6/ins[137] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[138]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[139] ),
    .A(\tapped_ring.c6/ins[138] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[139]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[140] ),
    .A(\tapped_ring.c6/ins[139] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[13]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[14] ),
    .A(\tapped_ring.c6/ins[13] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[140]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[141] ),
    .A(\tapped_ring.c6/ins[140] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[141]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[142] ),
    .A(\tapped_ring.c6/ins[141] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[142]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[143] ),
    .A(\tapped_ring.c6/ins[142] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[143]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[144] ),
    .A(\tapped_ring.c6/ins[143] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[144]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[145] ),
    .A(\tapped_ring.c6/ins[144] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[145]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[146] ),
    .A(\tapped_ring.c6/ins[145] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[146]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[147] ),
    .A(\tapped_ring.c6/ins[146] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[147]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[148] ),
    .A(\tapped_ring.c6/ins[147] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[148]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[149] ),
    .A(\tapped_ring.c6/ins[148] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[149]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[150] ),
    .A(\tapped_ring.c6/ins[149] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[14]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[15] ),
    .A(\tapped_ring.c6/ins[14] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[150]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[151] ),
    .A(\tapped_ring.c6/ins[150] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[151]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[152] ),
    .A(\tapped_ring.c6/ins[151] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[152]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[153] ),
    .A(\tapped_ring.c6/ins[152] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[153]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[154] ),
    .A(\tapped_ring.c6/ins[153] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[154]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[155] ),
    .A(\tapped_ring.c6/ins[154] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[155]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[156] ),
    .A(\tapped_ring.c6/ins[155] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[156]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[157] ),
    .A(\tapped_ring.c6/ins[156] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[157]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[158] ),
    .A(\tapped_ring.c6/ins[157] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[158]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[159] ),
    .A(\tapped_ring.c6/ins[158] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[159]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[160] ),
    .A(\tapped_ring.c6/ins[159] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[15]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[16] ),
    .A(\tapped_ring.c6/ins[15] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[160]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[161] ),
    .A(\tapped_ring.c6/ins[160] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[161]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[162] ),
    .A(\tapped_ring.c6/ins[161] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[162]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[163] ),
    .A(\tapped_ring.c6/ins[162] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[163]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[164] ),
    .A(\tapped_ring.c6/ins[163] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[164]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[165] ),
    .A(\tapped_ring.c6/ins[164] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[165]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[166] ),
    .A(\tapped_ring.c6/ins[165] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[166]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[167] ),
    .A(\tapped_ring.c6/ins[166] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[167]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[168] ),
    .A(\tapped_ring.c6/ins[167] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[168]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[169] ),
    .A(\tapped_ring.c6/ins[168] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[169]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[170] ),
    .A(\tapped_ring.c6/ins[169] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[16]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[17] ),
    .A(\tapped_ring.c6/ins[16] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[170]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[171] ),
    .A(\tapped_ring.c6/ins[170] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[171]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[172] ),
    .A(\tapped_ring.c6/ins[171] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[172]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[173] ),
    .A(\tapped_ring.c6/ins[172] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[173]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[174] ),
    .A(\tapped_ring.c6/ins[173] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[174]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[175] ),
    .A(\tapped_ring.c6/ins[174] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[175]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[176] ),
    .A(\tapped_ring.c6/ins[175] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[176]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[177] ),
    .A(\tapped_ring.c6/ins[176] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[177]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[178] ),
    .A(\tapped_ring.c6/ins[177] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[178]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[179] ),
    .A(\tapped_ring.c6/ins[178] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[179]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[180] ),
    .A(\tapped_ring.c6/ins[179] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[17]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[18] ),
    .A(\tapped_ring.c6/ins[17] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[180]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[181] ),
    .A(\tapped_ring.c6/ins[180] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[181]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[182] ),
    .A(\tapped_ring.c6/ins[181] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[182]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[183] ),
    .A(\tapped_ring.c6/ins[182] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[183]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[184] ),
    .A(\tapped_ring.c6/ins[183] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[184]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[185] ),
    .A(\tapped_ring.c6/ins[184] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[185]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[186] ),
    .A(\tapped_ring.c6/ins[185] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[186]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[187] ),
    .A(\tapped_ring.c6/ins[186] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[187]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[188] ),
    .A(\tapped_ring.c6/ins[187] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[188]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[189] ),
    .A(\tapped_ring.c6/ins[188] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[189]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[190] ),
    .A(\tapped_ring.c6/ins[189] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[18]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[19] ),
    .A(\tapped_ring.c6/ins[18] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[190]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[191] ),
    .A(\tapped_ring.c6/ins[190] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[191]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[192] ),
    .A(\tapped_ring.c6/ins[191] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[192]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[193] ),
    .A(\tapped_ring.c6/ins[192] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[193]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[194] ),
    .A(\tapped_ring.c6/ins[193] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[194]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[195] ),
    .A(\tapped_ring.c6/ins[194] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[195]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[196] ),
    .A(\tapped_ring.c6/ins[195] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[196]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[197] ),
    .A(\tapped_ring.c6/ins[196] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[197]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[198] ),
    .A(\tapped_ring.c6/ins[197] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[198]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[199] ),
    .A(\tapped_ring.c6/ins[198] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[199]/sky_inverter/_0_  (.Y(\tapped_ring.b301 ),
    .A(\tapped_ring.c6/ins[199] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[19]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[20] ),
    .A(\tapped_ring.c6/ins[19] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[2] ),
    .A(\tapped_ring.c6/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[20]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[21] ),
    .A(\tapped_ring.c6/ins[20] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[21]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[22] ),
    .A(\tapped_ring.c6/ins[21] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[22]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[23] ),
    .A(\tapped_ring.c6/ins[22] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[23]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[24] ),
    .A(\tapped_ring.c6/ins[23] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[24]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[25] ),
    .A(\tapped_ring.c6/ins[24] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[25]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[26] ),
    .A(\tapped_ring.c6/ins[25] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[26]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[27] ),
    .A(\tapped_ring.c6/ins[26] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[27]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[28] ),
    .A(\tapped_ring.c6/ins[27] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[28]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[29] ),
    .A(\tapped_ring.c6/ins[28] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[29]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[30] ),
    .A(\tapped_ring.c6/ins[29] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[3] ),
    .A(\tapped_ring.c6/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[30]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[31] ),
    .A(\tapped_ring.c6/ins[30] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[31]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[32] ),
    .A(\tapped_ring.c6/ins[31] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[32]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[33] ),
    .A(\tapped_ring.c6/ins[32] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[33]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[34] ),
    .A(\tapped_ring.c6/ins[33] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[34]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[35] ),
    .A(\tapped_ring.c6/ins[34] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[35]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[36] ),
    .A(\tapped_ring.c6/ins[35] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[36]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[37] ),
    .A(\tapped_ring.c6/ins[36] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[37]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[38] ),
    .A(\tapped_ring.c6/ins[37] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[38]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[39] ),
    .A(\tapped_ring.c6/ins[38] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[39]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[40] ),
    .A(\tapped_ring.c6/ins[39] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[4] ),
    .A(\tapped_ring.c6/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[40]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[41] ),
    .A(\tapped_ring.c6/ins[40] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[41]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[42] ),
    .A(\tapped_ring.c6/ins[41] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[42]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[43] ),
    .A(\tapped_ring.c6/ins[42] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[43]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[44] ),
    .A(\tapped_ring.c6/ins[43] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[44]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[45] ),
    .A(\tapped_ring.c6/ins[44] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[45]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[46] ),
    .A(\tapped_ring.c6/ins[45] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[46]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[47] ),
    .A(\tapped_ring.c6/ins[46] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[47]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[48] ),
    .A(\tapped_ring.c6/ins[47] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[48]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[49] ),
    .A(\tapped_ring.c6/ins[48] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[49]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[50] ),
    .A(\tapped_ring.c6/ins[49] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[5] ),
    .A(\tapped_ring.c6/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[50]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[51] ),
    .A(\tapped_ring.c6/ins[50] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[51]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[52] ),
    .A(\tapped_ring.c6/ins[51] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[52]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[53] ),
    .A(\tapped_ring.c6/ins[52] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[53]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[54] ),
    .A(\tapped_ring.c6/ins[53] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[54]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[55] ),
    .A(\tapped_ring.c6/ins[54] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[55]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[56] ),
    .A(\tapped_ring.c6/ins[55] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[56]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[57] ),
    .A(\tapped_ring.c6/ins[56] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[57]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[58] ),
    .A(\tapped_ring.c6/ins[57] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[58]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[59] ),
    .A(\tapped_ring.c6/ins[58] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[59]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[60] ),
    .A(\tapped_ring.c6/ins[59] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[6] ),
    .A(\tapped_ring.c6/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[60]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[61] ),
    .A(\tapped_ring.c6/ins[60] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[61]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[62] ),
    .A(\tapped_ring.c6/ins[61] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[62]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[63] ),
    .A(\tapped_ring.c6/ins[62] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[63]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[64] ),
    .A(\tapped_ring.c6/ins[63] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[64]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[65] ),
    .A(\tapped_ring.c6/ins[64] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[65]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[66] ),
    .A(\tapped_ring.c6/ins[65] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[66]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[67] ),
    .A(\tapped_ring.c6/ins[66] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[67]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[68] ),
    .A(\tapped_ring.c6/ins[67] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[68]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[69] ),
    .A(\tapped_ring.c6/ins[68] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[69]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[70] ),
    .A(\tapped_ring.c6/ins[69] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[7] ),
    .A(\tapped_ring.c6/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[70]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[71] ),
    .A(\tapped_ring.c6/ins[70] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[71]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[72] ),
    .A(\tapped_ring.c6/ins[71] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[72]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[73] ),
    .A(\tapped_ring.c6/ins[72] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[73]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[74] ),
    .A(\tapped_ring.c6/ins[73] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[74]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[75] ),
    .A(\tapped_ring.c6/ins[74] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[75]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[76] ),
    .A(\tapped_ring.c6/ins[75] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[76]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[77] ),
    .A(\tapped_ring.c6/ins[76] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[77]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[78] ),
    .A(\tapped_ring.c6/ins[77] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[78]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[79] ),
    .A(\tapped_ring.c6/ins[78] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[79]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[80] ),
    .A(\tapped_ring.c6/ins[79] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[8] ),
    .A(\tapped_ring.c6/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[80]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[81] ),
    .A(\tapped_ring.c6/ins[80] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[81]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[82] ),
    .A(\tapped_ring.c6/ins[81] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[82]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[83] ),
    .A(\tapped_ring.c6/ins[82] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[83]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[84] ),
    .A(\tapped_ring.c6/ins[83] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[84]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[85] ),
    .A(\tapped_ring.c6/ins[84] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[85]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[86] ),
    .A(\tapped_ring.c6/ins[85] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[86]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[87] ),
    .A(\tapped_ring.c6/ins[86] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[87]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[88] ),
    .A(\tapped_ring.c6/ins[87] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[88]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[89] ),
    .A(\tapped_ring.c6/ins[88] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[89]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[90] ),
    .A(\tapped_ring.c6/ins[89] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[9] ),
    .A(\tapped_ring.c6/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[90]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[91] ),
    .A(\tapped_ring.c6/ins[90] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[91]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[92] ),
    .A(\tapped_ring.c6/ins[91] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[92]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[93] ),
    .A(\tapped_ring.c6/ins[92] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[93]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[94] ),
    .A(\tapped_ring.c6/ins[93] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[94]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[95] ),
    .A(\tapped_ring.c6/ins[94] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[95]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[96] ),
    .A(\tapped_ring.c6/ins[95] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[96]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[97] ),
    .A(\tapped_ring.c6/ins[96] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[97]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[98] ),
    .A(\tapped_ring.c6/ins[97] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[98]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[99] ),
    .A(\tapped_ring.c6/ins[98] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[99]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[100] ),
    .A(\tapped_ring.c6/ins[99] ));
 sg13g2_inv_1 \tapped_ring.c6/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.c6/ins[10] ),
    .A(\tapped_ring.c6/ins[9] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[0]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[1] ),
    .A(\tapped_ring.b301 ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[100]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[101] ),
    .A(\tapped_ring.c7/ins[100] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[101]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[102] ),
    .A(\tapped_ring.c7/ins[101] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[102]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[103] ),
    .A(\tapped_ring.c7/ins[102] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[103]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[104] ),
    .A(\tapped_ring.c7/ins[103] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[104]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[105] ),
    .A(\tapped_ring.c7/ins[104] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[105]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[106] ),
    .A(\tapped_ring.c7/ins[105] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[106]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[107] ),
    .A(\tapped_ring.c7/ins[106] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[107]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[108] ),
    .A(\tapped_ring.c7/ins[107] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[108]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[109] ),
    .A(\tapped_ring.c7/ins[108] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[109]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[110] ),
    .A(\tapped_ring.c7/ins[109] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[10]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[11] ),
    .A(\tapped_ring.c7/ins[10] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[110]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[111] ),
    .A(\tapped_ring.c7/ins[110] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[111]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[112] ),
    .A(\tapped_ring.c7/ins[111] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[112]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[113] ),
    .A(\tapped_ring.c7/ins[112] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[113]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[114] ),
    .A(\tapped_ring.c7/ins[113] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[114]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[115] ),
    .A(\tapped_ring.c7/ins[114] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[115]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[116] ),
    .A(\tapped_ring.c7/ins[115] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[116]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[117] ),
    .A(\tapped_ring.c7/ins[116] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[117]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[118] ),
    .A(\tapped_ring.c7/ins[117] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[118]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[119] ),
    .A(\tapped_ring.c7/ins[118] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[119]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[120] ),
    .A(\tapped_ring.c7/ins[119] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[11]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[12] ),
    .A(\tapped_ring.c7/ins[11] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[120]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[121] ),
    .A(\tapped_ring.c7/ins[120] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[121]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[122] ),
    .A(\tapped_ring.c7/ins[121] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[122]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[123] ),
    .A(\tapped_ring.c7/ins[122] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[123]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[124] ),
    .A(\tapped_ring.c7/ins[123] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[124]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[125] ),
    .A(\tapped_ring.c7/ins[124] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[125]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[126] ),
    .A(\tapped_ring.c7/ins[125] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[126]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[127] ),
    .A(\tapped_ring.c7/ins[126] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[127]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[128] ),
    .A(\tapped_ring.c7/ins[127] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[128]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[129] ),
    .A(\tapped_ring.c7/ins[128] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[129]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[130] ),
    .A(\tapped_ring.c7/ins[129] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[12]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[13] ),
    .A(\tapped_ring.c7/ins[12] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[130]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[131] ),
    .A(\tapped_ring.c7/ins[130] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[131]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[132] ),
    .A(\tapped_ring.c7/ins[131] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[132]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[133] ),
    .A(\tapped_ring.c7/ins[132] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[133]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[134] ),
    .A(\tapped_ring.c7/ins[133] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[134]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[135] ),
    .A(\tapped_ring.c7/ins[134] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[135]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[136] ),
    .A(\tapped_ring.c7/ins[135] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[136]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[137] ),
    .A(\tapped_ring.c7/ins[136] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[137]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[138] ),
    .A(\tapped_ring.c7/ins[137] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[138]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[139] ),
    .A(\tapped_ring.c7/ins[138] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[139]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[140] ),
    .A(\tapped_ring.c7/ins[139] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[13]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[14] ),
    .A(\tapped_ring.c7/ins[13] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[140]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[141] ),
    .A(\tapped_ring.c7/ins[140] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[141]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[142] ),
    .A(\tapped_ring.c7/ins[141] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[142]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[143] ),
    .A(\tapped_ring.c7/ins[142] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[143]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[144] ),
    .A(\tapped_ring.c7/ins[143] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[144]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[145] ),
    .A(\tapped_ring.c7/ins[144] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[145]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[146] ),
    .A(\tapped_ring.c7/ins[145] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[146]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[147] ),
    .A(\tapped_ring.c7/ins[146] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[147]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[148] ),
    .A(\tapped_ring.c7/ins[147] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[148]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[149] ),
    .A(\tapped_ring.c7/ins[148] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[149]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[150] ),
    .A(\tapped_ring.c7/ins[149] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[14]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[15] ),
    .A(\tapped_ring.c7/ins[14] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[150]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[151] ),
    .A(\tapped_ring.c7/ins[150] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[151]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[152] ),
    .A(\tapped_ring.c7/ins[151] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[152]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[153] ),
    .A(\tapped_ring.c7/ins[152] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[153]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[154] ),
    .A(\tapped_ring.c7/ins[153] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[154]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[155] ),
    .A(\tapped_ring.c7/ins[154] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[155]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[156] ),
    .A(\tapped_ring.c7/ins[155] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[156]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[157] ),
    .A(\tapped_ring.c7/ins[156] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[157]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[158] ),
    .A(\tapped_ring.c7/ins[157] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[158]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[159] ),
    .A(\tapped_ring.c7/ins[158] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[159]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[160] ),
    .A(\tapped_ring.c7/ins[159] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[15]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[16] ),
    .A(\tapped_ring.c7/ins[15] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[160]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[161] ),
    .A(\tapped_ring.c7/ins[160] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[161]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[162] ),
    .A(\tapped_ring.c7/ins[161] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[162]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[163] ),
    .A(\tapped_ring.c7/ins[162] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[163]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[164] ),
    .A(\tapped_ring.c7/ins[163] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[164]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[165] ),
    .A(\tapped_ring.c7/ins[164] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[165]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[166] ),
    .A(\tapped_ring.c7/ins[165] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[166]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[167] ),
    .A(\tapped_ring.c7/ins[166] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[167]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[168] ),
    .A(\tapped_ring.c7/ins[167] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[168]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[169] ),
    .A(\tapped_ring.c7/ins[168] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[169]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[170] ),
    .A(\tapped_ring.c7/ins[169] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[16]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[17] ),
    .A(\tapped_ring.c7/ins[16] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[170]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[171] ),
    .A(\tapped_ring.c7/ins[170] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[171]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[172] ),
    .A(\tapped_ring.c7/ins[171] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[172]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[173] ),
    .A(\tapped_ring.c7/ins[172] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[173]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[174] ),
    .A(\tapped_ring.c7/ins[173] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[174]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[175] ),
    .A(\tapped_ring.c7/ins[174] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[175]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[176] ),
    .A(\tapped_ring.c7/ins[175] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[176]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[177] ),
    .A(\tapped_ring.c7/ins[176] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[177]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[178] ),
    .A(\tapped_ring.c7/ins[177] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[178]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[179] ),
    .A(\tapped_ring.c7/ins[178] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[179]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[180] ),
    .A(\tapped_ring.c7/ins[179] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[17]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[18] ),
    .A(\tapped_ring.c7/ins[17] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[180]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[181] ),
    .A(\tapped_ring.c7/ins[180] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[181]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[182] ),
    .A(\tapped_ring.c7/ins[181] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[182]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[183] ),
    .A(\tapped_ring.c7/ins[182] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[183]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[184] ),
    .A(\tapped_ring.c7/ins[183] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[184]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[185] ),
    .A(\tapped_ring.c7/ins[184] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[185]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[186] ),
    .A(\tapped_ring.c7/ins[185] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[186]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[187] ),
    .A(\tapped_ring.c7/ins[186] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[187]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[188] ),
    .A(\tapped_ring.c7/ins[187] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[188]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[189] ),
    .A(\tapped_ring.c7/ins[188] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[189]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[190] ),
    .A(\tapped_ring.c7/ins[189] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[18]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[19] ),
    .A(\tapped_ring.c7/ins[18] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[190]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[191] ),
    .A(\tapped_ring.c7/ins[190] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[191]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[192] ),
    .A(\tapped_ring.c7/ins[191] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[192]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[193] ),
    .A(\tapped_ring.c7/ins[192] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[193]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[194] ),
    .A(\tapped_ring.c7/ins[193] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[194]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[195] ),
    .A(\tapped_ring.c7/ins[194] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[195]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[196] ),
    .A(\tapped_ring.c7/ins[195] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[196]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[197] ),
    .A(\tapped_ring.c7/ins[196] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[197]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[198] ),
    .A(\tapped_ring.c7/ins[197] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[198]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[199] ),
    .A(\tapped_ring.c7/ins[198] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[199]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[200] ),
    .A(\tapped_ring.c7/ins[199] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[19]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[20] ),
    .A(\tapped_ring.c7/ins[19] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[1]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[2] ),
    .A(\tapped_ring.c7/ins[1] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[200]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[201] ),
    .A(\tapped_ring.c7/ins[200] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[201]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[202] ),
    .A(\tapped_ring.c7/ins[201] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[202]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[203] ),
    .A(\tapped_ring.c7/ins[202] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[203]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[204] ),
    .A(\tapped_ring.c7/ins[203] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[204]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[205] ),
    .A(\tapped_ring.c7/ins[204] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[205]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[206] ),
    .A(\tapped_ring.c7/ins[205] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[206]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[207] ),
    .A(\tapped_ring.c7/ins[206] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[207]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[208] ),
    .A(\tapped_ring.c7/ins[207] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[208]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[209] ),
    .A(\tapped_ring.c7/ins[208] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[209]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[210] ),
    .A(\tapped_ring.c7/ins[209] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[20]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[21] ),
    .A(\tapped_ring.c7/ins[20] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[210]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[211] ),
    .A(\tapped_ring.c7/ins[210] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[211]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[212] ),
    .A(\tapped_ring.c7/ins[211] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[212]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[213] ),
    .A(\tapped_ring.c7/ins[212] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[213]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[214] ),
    .A(\tapped_ring.c7/ins[213] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[214]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[215] ),
    .A(\tapped_ring.c7/ins[214] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[215]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[216] ),
    .A(\tapped_ring.c7/ins[215] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[216]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[217] ),
    .A(\tapped_ring.c7/ins[216] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[217]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[218] ),
    .A(\tapped_ring.c7/ins[217] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[218]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[219] ),
    .A(\tapped_ring.c7/ins[218] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[219]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[220] ),
    .A(\tapped_ring.c7/ins[219] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[21]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[22] ),
    .A(\tapped_ring.c7/ins[21] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[220]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[221] ),
    .A(\tapped_ring.c7/ins[220] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[221]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[222] ),
    .A(\tapped_ring.c7/ins[221] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[222]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[223] ),
    .A(\tapped_ring.c7/ins[222] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[223]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[224] ),
    .A(\tapped_ring.c7/ins[223] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[224]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[225] ),
    .A(\tapped_ring.c7/ins[224] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[225]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[226] ),
    .A(\tapped_ring.c7/ins[225] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[226]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[227] ),
    .A(\tapped_ring.c7/ins[226] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[227]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[228] ),
    .A(\tapped_ring.c7/ins[227] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[228]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[229] ),
    .A(\tapped_ring.c7/ins[228] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[229]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[230] ),
    .A(\tapped_ring.c7/ins[229] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[22]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[23] ),
    .A(\tapped_ring.c7/ins[22] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[230]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[231] ),
    .A(\tapped_ring.c7/ins[230] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[231]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[232] ),
    .A(\tapped_ring.c7/ins[231] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[232]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[233] ),
    .A(\tapped_ring.c7/ins[232] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[233]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[234] ),
    .A(\tapped_ring.c7/ins[233] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[234]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[235] ),
    .A(\tapped_ring.c7/ins[234] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[235]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[236] ),
    .A(\tapped_ring.c7/ins[235] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[236]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[237] ),
    .A(\tapped_ring.c7/ins[236] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[237]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[238] ),
    .A(\tapped_ring.c7/ins[237] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[238]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[239] ),
    .A(\tapped_ring.c7/ins[238] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[239]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[240] ),
    .A(\tapped_ring.c7/ins[239] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[23]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[24] ),
    .A(\tapped_ring.c7/ins[23] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[240]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[241] ),
    .A(\tapped_ring.c7/ins[240] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[241]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[242] ),
    .A(\tapped_ring.c7/ins[241] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[242]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[243] ),
    .A(\tapped_ring.c7/ins[242] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[243]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[244] ),
    .A(\tapped_ring.c7/ins[243] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[244]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[245] ),
    .A(\tapped_ring.c7/ins[244] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[245]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[246] ),
    .A(\tapped_ring.c7/ins[245] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[246]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[247] ),
    .A(\tapped_ring.c7/ins[246] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[247]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[248] ),
    .A(\tapped_ring.c7/ins[247] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[248]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[249] ),
    .A(\tapped_ring.c7/ins[248] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[249]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[250] ),
    .A(\tapped_ring.c7/ins[249] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[24]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[25] ),
    .A(\tapped_ring.c7/ins[24] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[250]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[251] ),
    .A(\tapped_ring.c7/ins[250] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[251]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[252] ),
    .A(\tapped_ring.c7/ins[251] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[252]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[253] ),
    .A(\tapped_ring.c7/ins[252] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[253]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[254] ),
    .A(\tapped_ring.c7/ins[253] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[254]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[255] ),
    .A(\tapped_ring.c7/ins[254] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[255]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[256] ),
    .A(\tapped_ring.c7/ins[255] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[256]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[257] ),
    .A(\tapped_ring.c7/ins[256] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[257]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[258] ),
    .A(\tapped_ring.c7/ins[257] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[258]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[259] ),
    .A(\tapped_ring.c7/ins[258] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[259]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[260] ),
    .A(\tapped_ring.c7/ins[259] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[25]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[26] ),
    .A(\tapped_ring.c7/ins[25] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[260]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[261] ),
    .A(\tapped_ring.c7/ins[260] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[261]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[262] ),
    .A(\tapped_ring.c7/ins[261] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[262]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[263] ),
    .A(\tapped_ring.c7/ins[262] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[263]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[264] ),
    .A(\tapped_ring.c7/ins[263] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[264]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[265] ),
    .A(\tapped_ring.c7/ins[264] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[265]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[266] ),
    .A(\tapped_ring.c7/ins[265] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[266]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[267] ),
    .A(\tapped_ring.c7/ins[266] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[267]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[268] ),
    .A(\tapped_ring.c7/ins[267] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[268]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[269] ),
    .A(\tapped_ring.c7/ins[268] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[269]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[270] ),
    .A(\tapped_ring.c7/ins[269] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[26]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[27] ),
    .A(\tapped_ring.c7/ins[26] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[270]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[271] ),
    .A(\tapped_ring.c7/ins[270] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[271]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[272] ),
    .A(\tapped_ring.c7/ins[271] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[272]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[273] ),
    .A(\tapped_ring.c7/ins[272] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[273]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[274] ),
    .A(\tapped_ring.c7/ins[273] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[274]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[275] ),
    .A(\tapped_ring.c7/ins[274] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[275]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[276] ),
    .A(\tapped_ring.c7/ins[275] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[276]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[277] ),
    .A(\tapped_ring.c7/ins[276] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[277]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[278] ),
    .A(\tapped_ring.c7/ins[277] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[278]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[279] ),
    .A(\tapped_ring.c7/ins[278] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[279]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[280] ),
    .A(\tapped_ring.c7/ins[279] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[27]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[28] ),
    .A(\tapped_ring.c7/ins[27] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[280]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[281] ),
    .A(\tapped_ring.c7/ins[280] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[281]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[282] ),
    .A(\tapped_ring.c7/ins[281] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[282]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[283] ),
    .A(\tapped_ring.c7/ins[282] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[283]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[284] ),
    .A(\tapped_ring.c7/ins[283] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[284]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[285] ),
    .A(\tapped_ring.c7/ins[284] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[285]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[286] ),
    .A(\tapped_ring.c7/ins[285] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[286]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[287] ),
    .A(\tapped_ring.c7/ins[286] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[287]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[288] ),
    .A(\tapped_ring.c7/ins[287] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[288]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[289] ),
    .A(\tapped_ring.c7/ins[288] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[289]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[290] ),
    .A(\tapped_ring.c7/ins[289] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[28]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[29] ),
    .A(\tapped_ring.c7/ins[28] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[290]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[291] ),
    .A(\tapped_ring.c7/ins[290] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[291]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[292] ),
    .A(\tapped_ring.c7/ins[291] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[292]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[293] ),
    .A(\tapped_ring.c7/ins[292] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[293]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[294] ),
    .A(\tapped_ring.c7/ins[293] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[294]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[295] ),
    .A(\tapped_ring.c7/ins[294] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[295]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[296] ),
    .A(\tapped_ring.c7/ins[295] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[296]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[297] ),
    .A(\tapped_ring.c7/ins[296] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[297]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[298] ),
    .A(\tapped_ring.c7/ins[297] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[298]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[299] ),
    .A(\tapped_ring.c7/ins[298] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[299]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[300] ),
    .A(\tapped_ring.c7/ins[299] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[29]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[30] ),
    .A(\tapped_ring.c7/ins[29] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[2]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[3] ),
    .A(\tapped_ring.c7/ins[2] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[300]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[301] ),
    .A(\tapped_ring.c7/ins[300] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[301]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[302] ),
    .A(\tapped_ring.c7/ins[301] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[302]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[303] ),
    .A(\tapped_ring.c7/ins[302] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[303]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[304] ),
    .A(\tapped_ring.c7/ins[303] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[304]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[305] ),
    .A(\tapped_ring.c7/ins[304] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[305]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[306] ),
    .A(\tapped_ring.c7/ins[305] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[306]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[307] ),
    .A(\tapped_ring.c7/ins[306] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[307]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[308] ),
    .A(\tapped_ring.c7/ins[307] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[308]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[309] ),
    .A(\tapped_ring.c7/ins[308] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[309]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[310] ),
    .A(\tapped_ring.c7/ins[309] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[30]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[31] ),
    .A(\tapped_ring.c7/ins[30] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[310]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[311] ),
    .A(\tapped_ring.c7/ins[310] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[311]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[312] ),
    .A(\tapped_ring.c7/ins[311] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[312]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[313] ),
    .A(\tapped_ring.c7/ins[312] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[313]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[314] ),
    .A(\tapped_ring.c7/ins[313] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[314]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[315] ),
    .A(\tapped_ring.c7/ins[314] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[315]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[316] ),
    .A(\tapped_ring.c7/ins[315] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[316]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[317] ),
    .A(\tapped_ring.c7/ins[316] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[317]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[318] ),
    .A(\tapped_ring.c7/ins[317] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[318]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[319] ),
    .A(\tapped_ring.c7/ins[318] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[319]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[320] ),
    .A(\tapped_ring.c7/ins[319] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[31]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[32] ),
    .A(\tapped_ring.c7/ins[31] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[320]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[321] ),
    .A(\tapped_ring.c7/ins[320] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[321]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[322] ),
    .A(\tapped_ring.c7/ins[321] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[322]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[323] ),
    .A(\tapped_ring.c7/ins[322] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[323]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[324] ),
    .A(\tapped_ring.c7/ins[323] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[324]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[325] ),
    .A(\tapped_ring.c7/ins[324] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[325]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[326] ),
    .A(\tapped_ring.c7/ins[325] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[326]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[327] ),
    .A(\tapped_ring.c7/ins[326] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[327]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[328] ),
    .A(\tapped_ring.c7/ins[327] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[328]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[329] ),
    .A(\tapped_ring.c7/ins[328] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[329]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[330] ),
    .A(\tapped_ring.c7/ins[329] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[32]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[33] ),
    .A(\tapped_ring.c7/ins[32] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[330]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[331] ),
    .A(\tapped_ring.c7/ins[330] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[331]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[332] ),
    .A(\tapped_ring.c7/ins[331] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[332]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[333] ),
    .A(\tapped_ring.c7/ins[332] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[333]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[334] ),
    .A(\tapped_ring.c7/ins[333] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[334]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[335] ),
    .A(\tapped_ring.c7/ins[334] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[335]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[336] ),
    .A(\tapped_ring.c7/ins[335] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[336]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[337] ),
    .A(\tapped_ring.c7/ins[336] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[337]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[338] ),
    .A(\tapped_ring.c7/ins[337] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[338]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[339] ),
    .A(\tapped_ring.c7/ins[338] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[339]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[340] ),
    .A(\tapped_ring.c7/ins[339] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[33]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[34] ),
    .A(\tapped_ring.c7/ins[33] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[340]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[341] ),
    .A(\tapped_ring.c7/ins[340] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[341]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[342] ),
    .A(\tapped_ring.c7/ins[341] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[342]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[343] ),
    .A(\tapped_ring.c7/ins[342] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[343]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[344] ),
    .A(\tapped_ring.c7/ins[343] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[344]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[345] ),
    .A(\tapped_ring.c7/ins[344] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[345]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[346] ),
    .A(\tapped_ring.c7/ins[345] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[346]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[347] ),
    .A(\tapped_ring.c7/ins[346] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[347]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[348] ),
    .A(\tapped_ring.c7/ins[347] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[348]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[349] ),
    .A(\tapped_ring.c7/ins[348] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[349]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[350] ),
    .A(\tapped_ring.c7/ins[349] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[34]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[35] ),
    .A(\tapped_ring.c7/ins[34] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[350]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[351] ),
    .A(\tapped_ring.c7/ins[350] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[351]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[352] ),
    .A(\tapped_ring.c7/ins[351] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[352]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[353] ),
    .A(\tapped_ring.c7/ins[352] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[353]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[354] ),
    .A(\tapped_ring.c7/ins[353] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[354]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[355] ),
    .A(\tapped_ring.c7/ins[354] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[355]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[356] ),
    .A(\tapped_ring.c7/ins[355] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[356]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[357] ),
    .A(\tapped_ring.c7/ins[356] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[357]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[358] ),
    .A(\tapped_ring.c7/ins[357] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[358]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[359] ),
    .A(\tapped_ring.c7/ins[358] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[359]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[360] ),
    .A(\tapped_ring.c7/ins[359] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[35]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[36] ),
    .A(\tapped_ring.c7/ins[35] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[360]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[361] ),
    .A(\tapped_ring.c7/ins[360] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[361]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[362] ),
    .A(\tapped_ring.c7/ins[361] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[362]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[363] ),
    .A(\tapped_ring.c7/ins[362] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[363]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[364] ),
    .A(\tapped_ring.c7/ins[363] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[364]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[365] ),
    .A(\tapped_ring.c7/ins[364] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[365]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[366] ),
    .A(\tapped_ring.c7/ins[365] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[366]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[367] ),
    .A(\tapped_ring.c7/ins[366] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[367]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[368] ),
    .A(\tapped_ring.c7/ins[367] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[368]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[369] ),
    .A(\tapped_ring.c7/ins[368] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[369]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[370] ),
    .A(\tapped_ring.c7/ins[369] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[36]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[37] ),
    .A(\tapped_ring.c7/ins[36] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[370]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[371] ),
    .A(\tapped_ring.c7/ins[370] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[371]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[372] ),
    .A(\tapped_ring.c7/ins[371] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[372]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[373] ),
    .A(\tapped_ring.c7/ins[372] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[373]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[374] ),
    .A(\tapped_ring.c7/ins[373] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[374]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[375] ),
    .A(\tapped_ring.c7/ins[374] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[375]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[376] ),
    .A(\tapped_ring.c7/ins[375] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[376]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[377] ),
    .A(\tapped_ring.c7/ins[376] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[377]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[378] ),
    .A(\tapped_ring.c7/ins[377] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[378]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[379] ),
    .A(\tapped_ring.c7/ins[378] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[379]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[380] ),
    .A(\tapped_ring.c7/ins[379] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[37]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[38] ),
    .A(\tapped_ring.c7/ins[37] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[380]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[381] ),
    .A(\tapped_ring.c7/ins[380] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[381]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[382] ),
    .A(\tapped_ring.c7/ins[381] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[382]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[383] ),
    .A(\tapped_ring.c7/ins[382] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[383]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[384] ),
    .A(\tapped_ring.c7/ins[383] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[384]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[385] ),
    .A(\tapped_ring.c7/ins[384] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[385]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[386] ),
    .A(\tapped_ring.c7/ins[385] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[386]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[387] ),
    .A(\tapped_ring.c7/ins[386] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[387]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[388] ),
    .A(\tapped_ring.c7/ins[387] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[388]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[389] ),
    .A(\tapped_ring.c7/ins[388] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[389]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[390] ),
    .A(\tapped_ring.c7/ins[389] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[38]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[39] ),
    .A(\tapped_ring.c7/ins[38] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[390]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[391] ),
    .A(\tapped_ring.c7/ins[390] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[391]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[392] ),
    .A(\tapped_ring.c7/ins[391] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[392]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[393] ),
    .A(\tapped_ring.c7/ins[392] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[393]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[394] ),
    .A(\tapped_ring.c7/ins[393] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[394]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[395] ),
    .A(\tapped_ring.c7/ins[394] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[395]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[396] ),
    .A(\tapped_ring.c7/ins[395] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[396]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[397] ),
    .A(\tapped_ring.c7/ins[396] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[397]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[398] ),
    .A(\tapped_ring.c7/ins[397] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[398]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[399] ),
    .A(\tapped_ring.c7/ins[398] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[399]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[400] ),
    .A(\tapped_ring.c7/ins[399] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[39]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[40] ),
    .A(\tapped_ring.c7/ins[39] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[3]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[4] ),
    .A(\tapped_ring.c7/ins[3] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[400]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[401] ),
    .A(\tapped_ring.c7/ins[400] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[401]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[402] ),
    .A(\tapped_ring.c7/ins[401] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[402]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[403] ),
    .A(\tapped_ring.c7/ins[402] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[403]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[404] ),
    .A(\tapped_ring.c7/ins[403] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[404]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[405] ),
    .A(\tapped_ring.c7/ins[404] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[405]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[406] ),
    .A(\tapped_ring.c7/ins[405] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[406]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[407] ),
    .A(\tapped_ring.c7/ins[406] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[407]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[408] ),
    .A(\tapped_ring.c7/ins[407] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[408]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[409] ),
    .A(\tapped_ring.c7/ins[408] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[409]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[410] ),
    .A(\tapped_ring.c7/ins[409] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[40]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[41] ),
    .A(\tapped_ring.c7/ins[40] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[410]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[411] ),
    .A(\tapped_ring.c7/ins[410] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[411]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[412] ),
    .A(\tapped_ring.c7/ins[411] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[412]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[413] ),
    .A(\tapped_ring.c7/ins[412] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[413]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[414] ),
    .A(\tapped_ring.c7/ins[413] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[414]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[415] ),
    .A(\tapped_ring.c7/ins[414] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[415]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[416] ),
    .A(\tapped_ring.c7/ins[415] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[416]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[417] ),
    .A(\tapped_ring.c7/ins[416] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[417]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[418] ),
    .A(\tapped_ring.c7/ins[417] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[418]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[419] ),
    .A(\tapped_ring.c7/ins[418] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[419]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[420] ),
    .A(\tapped_ring.c7/ins[419] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[41]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[42] ),
    .A(\tapped_ring.c7/ins[41] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[420]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[421] ),
    .A(\tapped_ring.c7/ins[420] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[421]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[422] ),
    .A(\tapped_ring.c7/ins[421] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[422]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[423] ),
    .A(\tapped_ring.c7/ins[422] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[423]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[424] ),
    .A(\tapped_ring.c7/ins[423] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[424]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[425] ),
    .A(\tapped_ring.c7/ins[424] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[425]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[426] ),
    .A(\tapped_ring.c7/ins[425] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[426]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[427] ),
    .A(\tapped_ring.c7/ins[426] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[427]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[428] ),
    .A(\tapped_ring.c7/ins[427] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[428]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[429] ),
    .A(\tapped_ring.c7/ins[428] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[429]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[430] ),
    .A(\tapped_ring.c7/ins[429] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[42]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[43] ),
    .A(\tapped_ring.c7/ins[42] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[430]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[431] ),
    .A(\tapped_ring.c7/ins[430] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[431]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[432] ),
    .A(\tapped_ring.c7/ins[431] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[432]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[433] ),
    .A(\tapped_ring.c7/ins[432] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[433]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[434] ),
    .A(\tapped_ring.c7/ins[433] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[434]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[435] ),
    .A(\tapped_ring.c7/ins[434] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[435]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[436] ),
    .A(\tapped_ring.c7/ins[435] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[436]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[437] ),
    .A(\tapped_ring.c7/ins[436] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[437]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[438] ),
    .A(\tapped_ring.c7/ins[437] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[438]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[439] ),
    .A(\tapped_ring.c7/ins[438] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[439]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[440] ),
    .A(\tapped_ring.c7/ins[439] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[43]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[44] ),
    .A(\tapped_ring.c7/ins[43] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[440]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[441] ),
    .A(\tapped_ring.c7/ins[440] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[441]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[442] ),
    .A(\tapped_ring.c7/ins[441] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[442]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[443] ),
    .A(\tapped_ring.c7/ins[442] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[443]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[444] ),
    .A(\tapped_ring.c7/ins[443] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[444]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[445] ),
    .A(\tapped_ring.c7/ins[444] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[445]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[446] ),
    .A(\tapped_ring.c7/ins[445] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[446]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[447] ),
    .A(\tapped_ring.c7/ins[446] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[447]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[448] ),
    .A(\tapped_ring.c7/ins[447] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[448]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[449] ),
    .A(\tapped_ring.c7/ins[448] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[449]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[450] ),
    .A(\tapped_ring.c7/ins[449] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[44]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[45] ),
    .A(\tapped_ring.c7/ins[44] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[450]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[451] ),
    .A(\tapped_ring.c7/ins[450] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[451]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[452] ),
    .A(\tapped_ring.c7/ins[451] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[452]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[453] ),
    .A(\tapped_ring.c7/ins[452] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[453]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[454] ),
    .A(\tapped_ring.c7/ins[453] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[454]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[455] ),
    .A(\tapped_ring.c7/ins[454] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[455]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[456] ),
    .A(\tapped_ring.c7/ins[455] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[456]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[457] ),
    .A(\tapped_ring.c7/ins[456] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[457]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[458] ),
    .A(\tapped_ring.c7/ins[457] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[458]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[459] ),
    .A(\tapped_ring.c7/ins[458] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[459]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[460] ),
    .A(\tapped_ring.c7/ins[459] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[45]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[46] ),
    .A(\tapped_ring.c7/ins[45] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[460]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[461] ),
    .A(\tapped_ring.c7/ins[460] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[461]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[462] ),
    .A(\tapped_ring.c7/ins[461] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[462]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[463] ),
    .A(\tapped_ring.c7/ins[462] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[463]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[464] ),
    .A(\tapped_ring.c7/ins[463] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[464]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[465] ),
    .A(\tapped_ring.c7/ins[464] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[465]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[466] ),
    .A(\tapped_ring.c7/ins[465] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[466]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[467] ),
    .A(\tapped_ring.c7/ins[466] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[467]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[468] ),
    .A(\tapped_ring.c7/ins[467] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[468]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[469] ),
    .A(\tapped_ring.c7/ins[468] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[469]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[470] ),
    .A(\tapped_ring.c7/ins[469] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[46]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[47] ),
    .A(\tapped_ring.c7/ins[46] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[470]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[471] ),
    .A(\tapped_ring.c7/ins[470] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[471]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[472] ),
    .A(\tapped_ring.c7/ins[471] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[472]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[473] ),
    .A(\tapped_ring.c7/ins[472] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[473]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[474] ),
    .A(\tapped_ring.c7/ins[473] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[474]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[475] ),
    .A(\tapped_ring.c7/ins[474] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[475]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[476] ),
    .A(\tapped_ring.c7/ins[475] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[476]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[477] ),
    .A(\tapped_ring.c7/ins[476] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[477]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[478] ),
    .A(\tapped_ring.c7/ins[477] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[478]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[479] ),
    .A(\tapped_ring.c7/ins[478] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[479]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[480] ),
    .A(\tapped_ring.c7/ins[479] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[47]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[48] ),
    .A(\tapped_ring.c7/ins[47] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[480]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[481] ),
    .A(\tapped_ring.c7/ins[480] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[481]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[482] ),
    .A(\tapped_ring.c7/ins[481] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[482]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[483] ),
    .A(\tapped_ring.c7/ins[482] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[483]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[484] ),
    .A(\tapped_ring.c7/ins[483] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[484]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[485] ),
    .A(\tapped_ring.c7/ins[484] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[485]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[486] ),
    .A(\tapped_ring.c7/ins[485] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[486]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[487] ),
    .A(\tapped_ring.c7/ins[486] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[487]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[488] ),
    .A(\tapped_ring.c7/ins[487] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[488]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[489] ),
    .A(\tapped_ring.c7/ins[488] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[489]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[490] ),
    .A(\tapped_ring.c7/ins[489] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[48]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[49] ),
    .A(\tapped_ring.c7/ins[48] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[490]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[491] ),
    .A(\tapped_ring.c7/ins[490] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[491]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[492] ),
    .A(\tapped_ring.c7/ins[491] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[492]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[493] ),
    .A(\tapped_ring.c7/ins[492] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[493]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[494] ),
    .A(\tapped_ring.c7/ins[493] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[494]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[495] ),
    .A(\tapped_ring.c7/ins[494] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[495]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[496] ),
    .A(\tapped_ring.c7/ins[495] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[496]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[497] ),
    .A(\tapped_ring.c7/ins[496] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[497]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[498] ),
    .A(\tapped_ring.c7/ins[497] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[498]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[499] ),
    .A(\tapped_ring.c7/ins[498] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[499]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[500] ),
    .A(\tapped_ring.c7/ins[499] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[49]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[50] ),
    .A(\tapped_ring.c7/ins[49] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[4]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[5] ),
    .A(\tapped_ring.c7/ins[4] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[500]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[501] ),
    .A(\tapped_ring.c7/ins[500] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[501]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[502] ),
    .A(\tapped_ring.c7/ins[501] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[502]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[503] ),
    .A(\tapped_ring.c7/ins[502] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[503]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[504] ),
    .A(\tapped_ring.c7/ins[503] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[504]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[505] ),
    .A(\tapped_ring.c7/ins[504] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[505]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[506] ),
    .A(\tapped_ring.c7/ins[505] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[506]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[507] ),
    .A(\tapped_ring.c7/ins[506] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[507]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[508] ),
    .A(\tapped_ring.c7/ins[507] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[508]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[509] ),
    .A(\tapped_ring.c7/ins[508] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[509]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[510] ),
    .A(\tapped_ring.c7/ins[509] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[50]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[51] ),
    .A(\tapped_ring.c7/ins[50] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[510]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[511] ),
    .A(\tapped_ring.c7/ins[510] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[511]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[512] ),
    .A(\tapped_ring.c7/ins[511] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[512]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[513] ),
    .A(\tapped_ring.c7/ins[512] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[513]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[514] ),
    .A(\tapped_ring.c7/ins[513] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[514]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[515] ),
    .A(\tapped_ring.c7/ins[514] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[515]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[516] ),
    .A(\tapped_ring.c7/ins[515] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[516]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[517] ),
    .A(\tapped_ring.c7/ins[516] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[517]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[518] ),
    .A(\tapped_ring.c7/ins[517] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[518]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[519] ),
    .A(\tapped_ring.c7/ins[518] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[519]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[520] ),
    .A(\tapped_ring.c7/ins[519] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[51]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[52] ),
    .A(\tapped_ring.c7/ins[51] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[520]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[521] ),
    .A(\tapped_ring.c7/ins[520] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[521]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[522] ),
    .A(\tapped_ring.c7/ins[521] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[522]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[523] ),
    .A(\tapped_ring.c7/ins[522] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[523]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[524] ),
    .A(\tapped_ring.c7/ins[523] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[524]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[525] ),
    .A(\tapped_ring.c7/ins[524] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[525]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[526] ),
    .A(\tapped_ring.c7/ins[525] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[526]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[527] ),
    .A(\tapped_ring.c7/ins[526] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[527]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[528] ),
    .A(\tapped_ring.c7/ins[527] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[528]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[529] ),
    .A(\tapped_ring.c7/ins[528] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[529]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[530] ),
    .A(\tapped_ring.c7/ins[529] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[52]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[53] ),
    .A(\tapped_ring.c7/ins[52] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[530]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[531] ),
    .A(\tapped_ring.c7/ins[530] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[531]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[532] ),
    .A(\tapped_ring.c7/ins[531] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[532]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[533] ),
    .A(\tapped_ring.c7/ins[532] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[533]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[534] ),
    .A(\tapped_ring.c7/ins[533] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[534]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[535] ),
    .A(\tapped_ring.c7/ins[534] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[535]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[536] ),
    .A(\tapped_ring.c7/ins[535] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[536]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[537] ),
    .A(\tapped_ring.c7/ins[536] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[537]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[538] ),
    .A(\tapped_ring.c7/ins[537] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[538]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[539] ),
    .A(\tapped_ring.c7/ins[538] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[539]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[540] ),
    .A(\tapped_ring.c7/ins[539] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[53]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[54] ),
    .A(\tapped_ring.c7/ins[53] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[540]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[541] ),
    .A(\tapped_ring.c7/ins[540] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[541]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[542] ),
    .A(\tapped_ring.c7/ins[541] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[542]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[543] ),
    .A(\tapped_ring.c7/ins[542] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[543]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[544] ),
    .A(\tapped_ring.c7/ins[543] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[544]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[545] ),
    .A(\tapped_ring.c7/ins[544] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[545]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[546] ),
    .A(\tapped_ring.c7/ins[545] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[546]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[547] ),
    .A(\tapped_ring.c7/ins[546] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[547]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[548] ),
    .A(\tapped_ring.c7/ins[547] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[548]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[549] ),
    .A(\tapped_ring.c7/ins[548] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[549]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[550] ),
    .A(\tapped_ring.c7/ins[549] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[54]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[55] ),
    .A(\tapped_ring.c7/ins[54] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[550]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[551] ),
    .A(\tapped_ring.c7/ins[550] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[551]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[552] ),
    .A(\tapped_ring.c7/ins[551] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[552]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[553] ),
    .A(\tapped_ring.c7/ins[552] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[553]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[554] ),
    .A(\tapped_ring.c7/ins[553] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[554]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[555] ),
    .A(\tapped_ring.c7/ins[554] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[555]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[556] ),
    .A(\tapped_ring.c7/ins[555] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[556]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[557] ),
    .A(\tapped_ring.c7/ins[556] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[557]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[558] ),
    .A(\tapped_ring.c7/ins[557] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[558]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[559] ),
    .A(\tapped_ring.c7/ins[558] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[559]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[560] ),
    .A(\tapped_ring.c7/ins[559] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[55]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[56] ),
    .A(\tapped_ring.c7/ins[55] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[560]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[561] ),
    .A(\tapped_ring.c7/ins[560] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[561]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[562] ),
    .A(\tapped_ring.c7/ins[561] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[562]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[563] ),
    .A(\tapped_ring.c7/ins[562] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[563]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[564] ),
    .A(\tapped_ring.c7/ins[563] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[564]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[565] ),
    .A(\tapped_ring.c7/ins[564] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[565]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[566] ),
    .A(\tapped_ring.c7/ins[565] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[566]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[567] ),
    .A(\tapped_ring.c7/ins[566] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[567]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[568] ),
    .A(\tapped_ring.c7/ins[567] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[568]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[569] ),
    .A(\tapped_ring.c7/ins[568] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[569]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[570] ),
    .A(\tapped_ring.c7/ins[569] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[56]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[57] ),
    .A(\tapped_ring.c7/ins[56] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[570]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[571] ),
    .A(\tapped_ring.c7/ins[570] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[571]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[572] ),
    .A(\tapped_ring.c7/ins[571] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[572]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[573] ),
    .A(\tapped_ring.c7/ins[572] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[573]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[574] ),
    .A(\tapped_ring.c7/ins[573] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[574]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[575] ),
    .A(\tapped_ring.c7/ins[574] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[575]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[576] ),
    .A(\tapped_ring.c7/ins[575] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[576]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[577] ),
    .A(\tapped_ring.c7/ins[576] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[577]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[578] ),
    .A(\tapped_ring.c7/ins[577] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[578]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[579] ),
    .A(\tapped_ring.c7/ins[578] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[579]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[580] ),
    .A(\tapped_ring.c7/ins[579] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[57]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[58] ),
    .A(\tapped_ring.c7/ins[57] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[580]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[581] ),
    .A(\tapped_ring.c7/ins[580] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[581]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[582] ),
    .A(\tapped_ring.c7/ins[581] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[582]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[583] ),
    .A(\tapped_ring.c7/ins[582] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[583]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[584] ),
    .A(\tapped_ring.c7/ins[583] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[584]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[585] ),
    .A(\tapped_ring.c7/ins[584] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[585]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[586] ),
    .A(\tapped_ring.c7/ins[585] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[586]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[587] ),
    .A(\tapped_ring.c7/ins[586] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[587]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[588] ),
    .A(\tapped_ring.c7/ins[587] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[588]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[589] ),
    .A(\tapped_ring.c7/ins[588] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[589]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[590] ),
    .A(\tapped_ring.c7/ins[589] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[58]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[59] ),
    .A(\tapped_ring.c7/ins[58] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[590]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[591] ),
    .A(\tapped_ring.c7/ins[590] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[591]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[592] ),
    .A(\tapped_ring.c7/ins[591] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[592]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[593] ),
    .A(\tapped_ring.c7/ins[592] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[593]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[594] ),
    .A(\tapped_ring.c7/ins[593] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[594]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[595] ),
    .A(\tapped_ring.c7/ins[594] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[595]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[596] ),
    .A(\tapped_ring.c7/ins[595] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[596]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[597] ),
    .A(\tapped_ring.c7/ins[596] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[597]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[598] ),
    .A(\tapped_ring.c7/ins[597] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[598]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[599] ),
    .A(\tapped_ring.c7/ins[598] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[599]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[600] ),
    .A(\tapped_ring.c7/ins[599] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[59]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[60] ),
    .A(\tapped_ring.c7/ins[59] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[5]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[6] ),
    .A(\tapped_ring.c7/ins[5] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[600]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[601] ),
    .A(\tapped_ring.c7/ins[600] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[601]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[602] ),
    .A(\tapped_ring.c7/ins[601] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[602]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[603] ),
    .A(\tapped_ring.c7/ins[602] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[603]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[604] ),
    .A(\tapped_ring.c7/ins[603] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[604]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[605] ),
    .A(\tapped_ring.c7/ins[604] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[605]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[606] ),
    .A(\tapped_ring.c7/ins[605] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[606]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[607] ),
    .A(\tapped_ring.c7/ins[606] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[607]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[608] ),
    .A(\tapped_ring.c7/ins[607] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[608]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[609] ),
    .A(\tapped_ring.c7/ins[608] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[609]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[610] ),
    .A(\tapped_ring.c7/ins[609] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[60]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[61] ),
    .A(\tapped_ring.c7/ins[60] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[610]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[611] ),
    .A(\tapped_ring.c7/ins[610] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[611]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[612] ),
    .A(\tapped_ring.c7/ins[611] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[612]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[613] ),
    .A(\tapped_ring.c7/ins[612] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[613]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[614] ),
    .A(\tapped_ring.c7/ins[613] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[614]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[615] ),
    .A(\tapped_ring.c7/ins[614] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[615]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[616] ),
    .A(\tapped_ring.c7/ins[615] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[616]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[617] ),
    .A(\tapped_ring.c7/ins[616] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[617]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[618] ),
    .A(\tapped_ring.c7/ins[617] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[618]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[619] ),
    .A(\tapped_ring.c7/ins[618] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[619]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[620] ),
    .A(\tapped_ring.c7/ins[619] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[61]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[62] ),
    .A(\tapped_ring.c7/ins[61] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[620]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[621] ),
    .A(\tapped_ring.c7/ins[620] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[621]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[622] ),
    .A(\tapped_ring.c7/ins[621] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[622]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[623] ),
    .A(\tapped_ring.c7/ins[622] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[623]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[624] ),
    .A(\tapped_ring.c7/ins[623] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[624]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[625] ),
    .A(\tapped_ring.c7/ins[624] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[625]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[626] ),
    .A(\tapped_ring.c7/ins[625] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[626]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[627] ),
    .A(\tapped_ring.c7/ins[626] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[627]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[628] ),
    .A(\tapped_ring.c7/ins[627] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[628]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[629] ),
    .A(\tapped_ring.c7/ins[628] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[629]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[630] ),
    .A(\tapped_ring.c7/ins[629] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[62]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[63] ),
    .A(\tapped_ring.c7/ins[62] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[630]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[631] ),
    .A(\tapped_ring.c7/ins[630] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[631]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[632] ),
    .A(\tapped_ring.c7/ins[631] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[632]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[633] ),
    .A(\tapped_ring.c7/ins[632] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[633]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[634] ),
    .A(\tapped_ring.c7/ins[633] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[634]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[635] ),
    .A(\tapped_ring.c7/ins[634] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[635]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[636] ),
    .A(\tapped_ring.c7/ins[635] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[636]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[637] ),
    .A(\tapped_ring.c7/ins[636] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[637]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[638] ),
    .A(\tapped_ring.c7/ins[637] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[638]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[639] ),
    .A(\tapped_ring.c7/ins[638] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[639]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[640] ),
    .A(\tapped_ring.c7/ins[639] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[63]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[64] ),
    .A(\tapped_ring.c7/ins[63] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[640]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[641] ),
    .A(\tapped_ring.c7/ins[640] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[641]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[642] ),
    .A(\tapped_ring.c7/ins[641] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[642]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[643] ),
    .A(\tapped_ring.c7/ins[642] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[643]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[644] ),
    .A(\tapped_ring.c7/ins[643] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[644]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[645] ),
    .A(\tapped_ring.c7/ins[644] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[645]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[646] ),
    .A(\tapped_ring.c7/ins[645] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[646]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[647] ),
    .A(\tapped_ring.c7/ins[646] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[647]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[648] ),
    .A(\tapped_ring.c7/ins[647] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[648]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[649] ),
    .A(\tapped_ring.c7/ins[648] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[649]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[650] ),
    .A(\tapped_ring.c7/ins[649] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[64]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[65] ),
    .A(\tapped_ring.c7/ins[64] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[650]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[651] ),
    .A(\tapped_ring.c7/ins[650] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[651]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[652] ),
    .A(\tapped_ring.c7/ins[651] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[652]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[653] ),
    .A(\tapped_ring.c7/ins[652] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[653]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[654] ),
    .A(\tapped_ring.c7/ins[653] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[654]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[655] ),
    .A(\tapped_ring.c7/ins[654] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[655]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[656] ),
    .A(\tapped_ring.c7/ins[655] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[656]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[657] ),
    .A(\tapped_ring.c7/ins[656] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[657]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[658] ),
    .A(\tapped_ring.c7/ins[657] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[658]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[659] ),
    .A(\tapped_ring.c7/ins[658] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[659]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[660] ),
    .A(\tapped_ring.c7/ins[659] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[65]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[66] ),
    .A(\tapped_ring.c7/ins[65] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[660]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[661] ),
    .A(\tapped_ring.c7/ins[660] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[661]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[662] ),
    .A(\tapped_ring.c7/ins[661] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[662]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[663] ),
    .A(\tapped_ring.c7/ins[662] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[663]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[664] ),
    .A(\tapped_ring.c7/ins[663] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[664]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[665] ),
    .A(\tapped_ring.c7/ins[664] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[665]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[666] ),
    .A(\tapped_ring.c7/ins[665] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[666]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[667] ),
    .A(\tapped_ring.c7/ins[666] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[667]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[668] ),
    .A(\tapped_ring.c7/ins[667] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[668]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[669] ),
    .A(\tapped_ring.c7/ins[668] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[669]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[670] ),
    .A(\tapped_ring.c7/ins[669] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[66]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[67] ),
    .A(\tapped_ring.c7/ins[66] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[670]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[671] ),
    .A(\tapped_ring.c7/ins[670] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[671]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[672] ),
    .A(\tapped_ring.c7/ins[671] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[672]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[673] ),
    .A(\tapped_ring.c7/ins[672] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[673]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[674] ),
    .A(\tapped_ring.c7/ins[673] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[674]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[675] ),
    .A(\tapped_ring.c7/ins[674] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[675]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[676] ),
    .A(\tapped_ring.c7/ins[675] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[676]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[677] ),
    .A(\tapped_ring.c7/ins[676] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[677]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[678] ),
    .A(\tapped_ring.c7/ins[677] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[678]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[679] ),
    .A(\tapped_ring.c7/ins[678] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[679]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[680] ),
    .A(\tapped_ring.c7/ins[679] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[67]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[68] ),
    .A(\tapped_ring.c7/ins[67] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[680]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[681] ),
    .A(\tapped_ring.c7/ins[680] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[681]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[682] ),
    .A(\tapped_ring.c7/ins[681] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[682]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[683] ),
    .A(\tapped_ring.c7/ins[682] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[683]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[684] ),
    .A(\tapped_ring.c7/ins[683] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[684]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[685] ),
    .A(\tapped_ring.c7/ins[684] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[685]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[686] ),
    .A(\tapped_ring.c7/ins[685] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[686]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[687] ),
    .A(\tapped_ring.c7/ins[686] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[687]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[688] ),
    .A(\tapped_ring.c7/ins[687] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[688]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[689] ),
    .A(\tapped_ring.c7/ins[688] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[689]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[690] ),
    .A(\tapped_ring.c7/ins[689] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[68]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[69] ),
    .A(\tapped_ring.c7/ins[68] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[690]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[691] ),
    .A(\tapped_ring.c7/ins[690] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[691]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[692] ),
    .A(\tapped_ring.c7/ins[691] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[692]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[693] ),
    .A(\tapped_ring.c7/ins[692] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[693]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[694] ),
    .A(\tapped_ring.c7/ins[693] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[694]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[695] ),
    .A(\tapped_ring.c7/ins[694] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[695]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[696] ),
    .A(\tapped_ring.c7/ins[695] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[696]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[697] ),
    .A(\tapped_ring.c7/ins[696] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[697]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[698] ),
    .A(\tapped_ring.c7/ins[697] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[698]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[699] ),
    .A(\tapped_ring.c7/ins[698] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[699]/sky_inverter/_0_  (.Y(\tapped_ring.b1001 ),
    .A(\tapped_ring.c7/ins[699] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[69]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[70] ),
    .A(\tapped_ring.c7/ins[69] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[6]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[7] ),
    .A(\tapped_ring.c7/ins[6] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[70]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[71] ),
    .A(\tapped_ring.c7/ins[70] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[71]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[72] ),
    .A(\tapped_ring.c7/ins[71] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[72]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[73] ),
    .A(\tapped_ring.c7/ins[72] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[73]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[74] ),
    .A(\tapped_ring.c7/ins[73] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[74]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[75] ),
    .A(\tapped_ring.c7/ins[74] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[75]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[76] ),
    .A(\tapped_ring.c7/ins[75] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[76]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[77] ),
    .A(\tapped_ring.c7/ins[76] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[77]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[78] ),
    .A(\tapped_ring.c7/ins[77] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[78]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[79] ),
    .A(\tapped_ring.c7/ins[78] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[79]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[80] ),
    .A(\tapped_ring.c7/ins[79] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[7]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[8] ),
    .A(\tapped_ring.c7/ins[7] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[80]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[81] ),
    .A(\tapped_ring.c7/ins[80] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[81]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[82] ),
    .A(\tapped_ring.c7/ins[81] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[82]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[83] ),
    .A(\tapped_ring.c7/ins[82] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[83]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[84] ),
    .A(\tapped_ring.c7/ins[83] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[84]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[85] ),
    .A(\tapped_ring.c7/ins[84] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[85]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[86] ),
    .A(\tapped_ring.c7/ins[85] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[86]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[87] ),
    .A(\tapped_ring.c7/ins[86] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[87]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[88] ),
    .A(\tapped_ring.c7/ins[87] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[88]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[89] ),
    .A(\tapped_ring.c7/ins[88] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[89]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[90] ),
    .A(\tapped_ring.c7/ins[89] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[8]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[9] ),
    .A(\tapped_ring.c7/ins[8] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[90]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[91] ),
    .A(\tapped_ring.c7/ins[90] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[91]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[92] ),
    .A(\tapped_ring.c7/ins[91] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[92]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[93] ),
    .A(\tapped_ring.c7/ins[92] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[93]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[94] ),
    .A(\tapped_ring.c7/ins[93] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[94]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[95] ),
    .A(\tapped_ring.c7/ins[94] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[95]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[96] ),
    .A(\tapped_ring.c7/ins[95] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[96]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[97] ),
    .A(\tapped_ring.c7/ins[96] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[97]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[98] ),
    .A(\tapped_ring.c7/ins[97] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[98]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[99] ),
    .A(\tapped_ring.c7/ins[98] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[99]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[100] ),
    .A(\tapped_ring.c7/ins[99] ));
 sg13g2_inv_1 \tapped_ring.c7/inv_array[9]/sky_inverter/_0_  (.Y(\tapped_ring.c7/ins[10] ),
    .A(\tapped_ring.c7/ins[9] ));
 sg13g2_inv_1 \tapped_ring.start/sky_inverter/_0_  (.Y(\tapped_ring.b1 ),
    .A(\tapped_ring.b0 ));
 sg13g2_buf_2 fanout1 (.A(osc),
    .X(net1));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net2));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net3));
 sg13g2_buf_2 input3 (.A(ui_in[0]),
    .X(net4));
 sg13g2_buf_1 input4 (.A(ui_in[1]),
    .X(net5));
 sg13g2_buf_2 input5 (.A(ui_in[2]),
    .X(net6));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net7));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net8));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net9));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net10));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net11));
 sg13g2_buf_1 input11 (.A(uio_in[0]),
    .X(net12));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net13));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net14));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net15));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net16));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net17));
 sg13g2_buf_1 input17 (.A(uio_in[6]),
    .X(net18));
 sg13g2_buf_1 input18 (.A(uio_in[7]),
    .X(net19));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc3_19 (.L_LO(net20));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_4 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_4 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_4 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_278 ();
 sg13g2_decap_8 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_decap_4 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_326 ();
 sg13g2_decap_4 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_4 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_4 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_4 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_4 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_271 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_4 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_8 FILLER_26_204 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_275 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_decap_8 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_decap_4 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_195 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_decap_4 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_4 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_decap_4 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_132 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_decap_4 FILLER_30_159 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_171 ();
 sg13g2_decap_8 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_4 FILLER_30_384 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_4 FILLER_31_281 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_4 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_4 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_decap_4 FILLER_32_234 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_279 ();
 sg13g2_decap_4 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_4 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_fill_1 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_87 ();
 sg13g2_decap_8 FILLER_33_94 ();
 sg13g2_decap_8 FILLER_33_101 ();
 sg13g2_fill_2 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_190 ();
 sg13g2_decap_8 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_decap_4 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_332 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_decap_4 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_128 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_decap_4 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_decap_4 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_4 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_319 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_4 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_169 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_1 FILLER_35_258 ();
 sg13g2_decap_4 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_decap_4 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_decap_8 FILLER_36_150 ();
 sg13g2_decap_4 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_decap_4 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_272 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_decap_4 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_351 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_125 ();
 sg13g2_decap_8 FILLER_37_132 ();
 sg13g2_decap_8 FILLER_37_139 ();
 sg13g2_decap_8 FILLER_37_146 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_160 ();
 sg13g2_decap_4 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net41;
 assign uio_oe[1] = net20;
 assign uio_oe[2] = net21;
 assign uio_oe[3] = net22;
 assign uio_oe[4] = net23;
 assign uio_oe[5] = net24;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net26;
 assign uio_out[1] = net27;
 assign uio_out[2] = net28;
 assign uio_out[3] = net29;
 assign uio_out[4] = net30;
 assign uio_out[5] = net31;
 assign uio_out[6] = net32;
 assign uio_out[7] = net33;
endmodule

module tt_um_daobaanh_rng (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \TRNG_inst.TX_Active ;
 wire \TRNG_inst.TX_Byte[0] ;
 wire \TRNG_inst.TX_Byte[1] ;
 wire \TRNG_inst.TX_Byte[2] ;
 wire \TRNG_inst.TX_Byte[3] ;
 wire \TRNG_inst.TX_Byte[4] ;
 wire \TRNG_inst.TX_Byte[5] ;
 wire \TRNG_inst.TX_Byte[6] ;
 wire \TRNG_inst.TX_Byte[7] ;
 wire \TRNG_inst.TX_DV ;
 wire \TRNG_inst.TX_Serial ;
 wire \TRNG_inst.U1_TRNG.i_rst ;
 wire \TRNG_inst.U1_TRNG.o_RNG ;
 wire \TRNG_inst.U1_TRNG.o_data[0] ;
 wire \TRNG_inst.U1_TRNG.o_data[10] ;
 wire \TRNG_inst.U1_TRNG.o_data[11] ;
 wire \TRNG_inst.U1_TRNG.o_data[12] ;
 wire \TRNG_inst.U1_TRNG.o_data[13] ;
 wire \TRNG_inst.U1_TRNG.o_data[14] ;
 wire \TRNG_inst.U1_TRNG.o_data[15] ;
 wire \TRNG_inst.U1_TRNG.o_data[16] ;
 wire \TRNG_inst.U1_TRNG.o_data[17] ;
 wire \TRNG_inst.U1_TRNG.o_data[18] ;
 wire \TRNG_inst.U1_TRNG.o_data[19] ;
 wire \TRNG_inst.U1_TRNG.o_data[1] ;
 wire \TRNG_inst.U1_TRNG.o_data[20] ;
 wire \TRNG_inst.U1_TRNG.o_data[21] ;
 wire \TRNG_inst.U1_TRNG.o_data[22] ;
 wire \TRNG_inst.U1_TRNG.o_data[23] ;
 wire \TRNG_inst.U1_TRNG.o_data[24] ;
 wire \TRNG_inst.U1_TRNG.o_data[25] ;
 wire \TRNG_inst.U1_TRNG.o_data[26] ;
 wire \TRNG_inst.U1_TRNG.o_data[27] ;
 wire \TRNG_inst.U1_TRNG.o_data[28] ;
 wire \TRNG_inst.U1_TRNG.o_data[29] ;
 wire \TRNG_inst.U1_TRNG.o_data[2] ;
 wire \TRNG_inst.U1_TRNG.o_data[30] ;
 wire \TRNG_inst.U1_TRNG.o_data[31] ;
 wire \TRNG_inst.U1_TRNG.o_data[3] ;
 wire \TRNG_inst.U1_TRNG.o_data[4] ;
 wire \TRNG_inst.U1_TRNG.o_data[5] ;
 wire \TRNG_inst.U1_TRNG.o_data[6] ;
 wire \TRNG_inst.U1_TRNG.o_data[7] ;
 wire \TRNG_inst.U1_TRNG.o_data[8] ;
 wire \TRNG_inst.U1_TRNG.o_data[9] ;
 wire \TRNG_inst.U1_TRNG.w[10] ;
 wire \TRNG_inst.U1_TRNG.w[1] ;
 wire \TRNG_inst.U1_TRNG.w[2] ;
 wire \TRNG_inst.U1_TRNG.w[3] ;
 wire \TRNG_inst.U1_TRNG.w[4] ;
 wire \TRNG_inst.U1_TRNG.w[5] ;
 wire \TRNG_inst.U1_TRNG.w[6] ;
 wire \TRNG_inst.U1_TRNG.w[7] ;
 wire \TRNG_inst.U1_TRNG.w[8] ;
 wire \TRNG_inst.U1_TRNG.w[9] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[2] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[0] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[3] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[4] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[6] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[7] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[8] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[0] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[1] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[2] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[3] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[4] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[5] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[6] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[7] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_DV ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_RX_Data_R ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[1] ;
 wire \TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[2] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[2] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[1] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[8] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[9] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[1] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[2] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[0] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[1] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[2] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[3] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[4] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[5] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[6] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[7] ;
 wire \TRNG_inst.U2_UART_interface.TX_part.r_TX_Done ;
 wire \TRNG_inst.U3_Main_controller.cnt_bytes[0] ;
 wire \TRNG_inst.U3_Main_controller.cnt_bytes[1] ;
 wire \TRNG_inst.U3_Main_controller.cnt_bytes[2] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[0] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[10] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[1] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[2] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[3] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[4] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[5] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[6] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[7] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[8] ;
 wire \TRNG_inst.U3_Main_controller.cnt_delay[9] ;
 wire \TRNG_inst.U3_Main_controller.led ;
 wire \TRNG_inst.U3_Main_controller.state[0] ;
 wire \TRNG_inst.U3_Main_controller.state[1] ;
 wire \TRNG_inst.U3_Main_controller.state[2] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[0] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[10] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[11] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[12] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[13] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[14] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[15] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[16] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[17] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[18] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[19] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[1] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[20] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[21] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[22] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[23] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[24] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[25] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[26] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[27] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[28] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[29] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[2] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[30] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[31] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[3] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[4] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[5] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[6] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[7] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[8] ;
 wire \TRNG_inst.U3_Main_controller.tmp_reg[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire clknet_0_clk;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[0] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[10] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[11] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[12] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[13] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[14] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[15] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[16] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[17] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[18] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[19] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[1] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[20] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[21] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[22] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[23] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[24] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[25] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[26] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[27] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[28] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[29] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[2] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[30] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[3] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[4] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[5] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[6] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[7] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[8] ;
 wire \TRNG_inst.U1_TRNG.RG_part/i_r[9] ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_1_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_0_ ;
 wire \TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_1_ ;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;

 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_00_  (.B(net206),
    .A(uo_out[1]),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[0] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_01_  (.B(net198),
    .A(\TRNG_inst.U1_TRNG.w[1] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[2] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_02_  (.B(net291),
    .A(\TRNG_inst.U1_TRNG.w[2] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[4] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_03_  (.B(net194),
    .A(\TRNG_inst.U1_TRNG.w[3] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[6] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_04_  (.B(net197),
    .A(\TRNG_inst.U1_TRNG.w[4] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[8] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_05_  (.B(net314),
    .A(\TRNG_inst.U1_TRNG.w[5] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[10] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_06_  (.B(net332),
    .A(\TRNG_inst.U1_TRNG.w[6] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[12] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_07_  (.B(net201),
    .A(\TRNG_inst.U1_TRNG.w[7] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[14] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_08_  (.B(net235),
    .A(\TRNG_inst.U1_TRNG.o_data[13] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[17] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_09_  (.B(net278),
    .A(\TRNG_inst.U1_TRNG.o_data[11] ),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[20] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_10_  (.B(net217),
    .A(net184),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[23] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_11_  (.B(net215),
    .A(net291),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[25] ));
 sg13g2_xor2_1 \TRNG_inst.U1_TRNG.RG_part/_12_  (.B(net199),
    .A(net185),
    .X(\TRNG_inst.U1_TRNG.RG_part/i_r[28] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_13_  (.A(net181),
    .X(\TRNG_inst.U1_TRNG.o_data[0] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_14_  (.A(net185),
    .X(\TRNG_inst.U1_TRNG.o_data[2] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_15_  (.A(net182),
    .X(\TRNG_inst.U1_TRNG.o_data[4] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_16_  (.A(net168),
    .X(\TRNG_inst.U1_TRNG.o_data[6] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_17_  (.A(net184),
    .X(\TRNG_inst.U1_TRNG.o_data[8] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_18_  (.A(net175),
    .X(\TRNG_inst.U1_TRNG.o_data[10] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_19_  (.A(net174),
    .X(\TRNG_inst.U1_TRNG.o_data[12] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_20_  (.A(net169),
    .X(\TRNG_inst.U1_TRNG.o_data[14] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_21_  (.A(net178),
    .X(\TRNG_inst.U1_TRNG.o_data[16] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_22_  (.A(net180),
    .X(\TRNG_inst.U1_TRNG.o_data[17] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_23_  (.A(net171),
    .X(\TRNG_inst.U1_TRNG.o_data[19] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_24_  (.A(net172),
    .X(\TRNG_inst.U1_TRNG.o_data[20] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_25_  (.A(net173),
    .X(\TRNG_inst.U1_TRNG.o_data[22] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_26_  (.A(net167),
    .X(\TRNG_inst.U1_TRNG.o_data[23] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_27_  (.A(net170),
    .X(\TRNG_inst.U1_TRNG.o_data[25] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_28_  (.A(net176),
    .X(\TRNG_inst.U1_TRNG.o_data[27] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_29_  (.A(net177),
    .X(\TRNG_inst.U1_TRNG.o_data[28] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_30_  (.A(net183),
    .X(\TRNG_inst.U1_TRNG.o_data[30] ));
 sg13g2_buf_1 \TRNG_inst.U1_TRNG.RG_part/_31_  (.A(net179),
    .X(\TRNG_inst.U1_TRNG.o_data[31] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_3_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[0] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[0].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_RNG ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_0_ ),
    .A(net116));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_3_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[10] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[10].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[9] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_3_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_0_ ),
    .D(net174),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[11].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[11] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_3_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[12] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[12].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[11] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_3_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_0_ ),
    .D(net169),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[13].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[13] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_3_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[14] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[14].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[13] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_3_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_0_ ),
    .D(net178),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[15].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[15] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_3_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_0_ ),
    .D(net180),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[16].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[15] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_3_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_0_ ),
    .D(net236),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[17].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[16] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_3_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_0_ ),
    .D(net171),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[18].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[18] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_3_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_0_ ),
    .D(net172),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[19].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[18] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_3_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_0_ ),
    .D(net185),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[1].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[1] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_3_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_0_ ),
    .D(net279),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[20].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[19] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_0_ ),
    .A(net116));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_3_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_0_ ),
    .D(net173),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[21].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[21] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_0_ ),
    .A(net116));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_3_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_0_ ),
    .D(net167),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[22].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[21] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_3_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[23] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[23].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[22] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_3_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_0_ ),
    .D(net170),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[24].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[24] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_0_ ),
    .A(net117));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_3_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[25] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[25].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[24] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_3_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_0_ ),
    .D(net176),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[26].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[26] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_3_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_0_ ),
    .D(net177),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[27].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[26] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_0_ ),
    .A(net119));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_3_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[28] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[28].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[27] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_0_ ),
    .A(net119));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_3_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_0_ ),
    .D(net183),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[29].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[29] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_3_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[2] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[2].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[1] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_0_ ),
    .A(net119));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_3_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_0_ ),
    .D(net179),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[30].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[29] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_3_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_0_ ),
    .D(net181),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[31].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[30] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_3_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_0_ ),
    .D(net182),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[3].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[3] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_0_ ),
    .A(net118));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_3_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[4] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[4].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[3] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_0_ ),
    .A(net120));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_3_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_0_ ),
    .D(net168),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[5].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[5] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_0_ ),
    .A(net120));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_3_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[6] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[6].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[5] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_0_ ),
    .A(net116));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_3_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_0_ ),
    .D(net184),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[7].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[7] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_3_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_0_ ),
    .D(\TRNG_inst.U1_TRNG.RG_part/i_r[8] ),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[8].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.RG_part/i_r[7] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_2_  (.Y(\TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_0_ ),
    .A(net115));
 sg13g2_dfrbp_1 \TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_3_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(\TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_0_ ),
    .D(net175),
    .Q_N(\TRNG_inst.U1_TRNG.RG_part/genblk1[9].FF/_1_ ),
    .Q(\TRNG_inst.U1_TRNG.o_data[9] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[0].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[1] ),
    .A(uo_out[1]));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[1].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[2] ),
    .A(\TRNG_inst.U1_TRNG.w[1] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[2].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[3] ),
    .A(\TRNG_inst.U1_TRNG.w[2] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[3].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[4] ),
    .A(\TRNG_inst.U1_TRNG.w[3] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[4].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[5] ),
    .A(\TRNG_inst.U1_TRNG.w[4] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[5].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[6] ),
    .A(\TRNG_inst.U1_TRNG.w[5] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[6].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[7] ),
    .A(\TRNG_inst.U1_TRNG.w[6] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[7].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[8] ),
    .A(\TRNG_inst.U1_TRNG.w[7] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[8].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[9] ),
    .A(\TRNG_inst.U1_TRNG.w[8] ));
 sg13g2_inv_1 \TRNG_inst.U1_TRNG.RO_part/genblk1[9].not1/_0_  (.Y(\TRNG_inst.U1_TRNG.w[10] ),
    .A(\TRNG_inst.U1_TRNG.w[9] ));
 sg13g2_nand2_2 \TRNG_inst.U1_TRNG.RO_part/nand1/_0_  (.Y(uo_out[1]),
    .A(net1),
    .B(\TRNG_inst.U1_TRNG.w[10] ));
 sg13g2_inv_1 _0678_ (.Y(_0127_),
    .A(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ));
 sg13g2_inv_1 _0679_ (.Y(_0128_),
    .A(net207));
 sg13g2_inv_1 _0680_ (.Y(_0129_),
    .A(net335));
 sg13g2_inv_1 _0681_ (.Y(_0130_),
    .A(\TRNG_inst.U3_Main_controller.state[0] ));
 sg13g2_inv_1 _0682_ (.Y(_0131_),
    .A(net347));
 sg13g2_inv_1 _0683_ (.Y(_0132_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ));
 sg13g2_inv_1 _0684_ (.Y(_0133_),
    .A(_0002_));
 sg13g2_inv_1 _0685_ (.Y(_0134_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ));
 sg13g2_inv_1 _0686_ (.Y(_0135_),
    .A(net111));
 sg13g2_inv_1 _0687_ (.Y(_0136_),
    .A(net302));
 sg13g2_inv_1 _0688_ (.Y(_0137_),
    .A(net379));
 sg13g2_inv_1 _0689_ (.Y(_0138_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ));
 sg13g2_inv_1 _0690_ (.Y(_0139_),
    .A(net345));
 sg13g2_inv_1 _0691_ (.Y(_0140_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ));
 sg13g2_inv_1 _0692_ (.Y(_0141_),
    .A(net330));
 sg13g2_inv_1 _0693_ (.Y(_0142_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ));
 sg13g2_inv_1 _0694_ (.Y(_0143_),
    .A(net204));
 sg13g2_inv_1 _0695_ (.Y(_0144_),
    .A(net315));
 sg13g2_inv_1 _0696_ (.Y(_0145_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ));
 sg13g2_inv_1 _0697_ (.Y(_0146_),
    .A(net222));
 sg13g2_inv_1 _0698_ (.Y(_0147_),
    .A(net202));
 sg13g2_inv_1 _0699_ (.Y(_0148_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[5] ));
 sg13g2_inv_1 _0700_ (.Y(_0149_),
    .A(\TRNG_inst.U3_Main_controller.tmp_reg[24] ));
 sg13g2_inv_1 _0701_ (.Y(_0150_),
    .A(net242));
 sg13g2_inv_1 _0702_ (.Y(_0151_),
    .A(net245));
 sg13g2_inv_1 _0703_ (.Y(_0152_),
    .A(net310));
 sg13g2_inv_1 _0704_ (.Y(_0153_),
    .A(net253));
 sg13g2_inv_1 _0705_ (.Y(_0154_),
    .A(net262));
 sg13g2_inv_1 _0706_ (.Y(_0155_),
    .A(net224));
 sg13g2_inv_1 _0707_ (.Y(_0156_),
    .A(net214));
 sg13g2_inv_1 _0708_ (.Y(_0157_),
    .A(\TRNG_inst.U3_Main_controller.tmp_reg[26] ));
 sg13g2_inv_1 _0709_ (.Y(_0158_),
    .A(net254));
 sg13g2_inv_1 _0710_ (.Y(_0159_),
    .A(net263));
 sg13g2_inv_1 _0711_ (.Y(_0160_),
    .A(net313));
 sg13g2_inv_1 _0712_ (.Y(_0161_),
    .A(net290));
 sg13g2_inv_1 _0713_ (.Y(_0162_),
    .A(net287));
 sg13g2_inv_1 _0714_ (.Y(_0163_),
    .A(net296));
 sg13g2_inv_1 _0715_ (.Y(_0164_),
    .A(net221));
 sg13g2_inv_1 _0716_ (.Y(_0165_),
    .A(net234));
 sg13g2_inv_1 _0717_ (.Y(_0166_),
    .A(net298));
 sg13g2_inv_1 _0718_ (.Y(_0167_),
    .A(net273));
 sg13g2_inv_1 _0719_ (.Y(_0168_),
    .A(net283));
 sg13g2_inv_1 _0720_ (.Y(_0169_),
    .A(net228));
 sg13g2_inv_1 _0721_ (.Y(_0170_),
    .A(net259));
 sg13g2_inv_1 _0722_ (.Y(_0171_),
    .A(net274));
 sg13g2_inv_1 _0723_ (.Y(_0172_),
    .A(net267));
 sg13g2_inv_1 _0724_ (.Y(_0173_),
    .A(net252));
 sg13g2_inv_1 _0725_ (.Y(_0174_),
    .A(net246));
 sg13g2_inv_1 _0726_ (.Y(_0175_),
    .A(net301));
 sg13g2_inv_1 _0727_ (.Y(_0176_),
    .A(net282));
 sg13g2_inv_1 _0728_ (.Y(_0177_),
    .A(net249));
 sg13g2_inv_1 _0729_ (.Y(_0178_),
    .A(net230));
 sg13g2_inv_1 _0730_ (.Y(_0179_),
    .A(net229));
 sg13g2_inv_1 _0731_ (.Y(_0180_),
    .A(net200));
 sg13g2_inv_1 _0732_ (.Y(_0181_),
    .A(net269));
 sg13g2_inv_1 _0733_ (.Y(_0182_),
    .A(net120));
 sg13g2_nand3b_1 _0734_ (.B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ),
    .C(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ),
    .Y(_0183_),
    .A_N(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ));
 sg13g2_or2_1 _0735_ (.X(_0184_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ),
    .A(net318));
 sg13g2_nor2b_1 _0736_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .B_N(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ),
    .Y(_0185_));
 sg13g2_nand2b_1 _0737_ (.Y(_0186_),
    .B(_0006_),
    .A_N(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ));
 sg13g2_a21oi_1 _0738_ (.A1(_0184_),
    .A2(_0185_),
    .Y(_0187_),
    .B1(_0186_));
 sg13g2_o21ai_1 _0739_ (.B1(net389),
    .Y(_0188_),
    .A1(_0183_),
    .A2(_0187_));
 sg13g2_and2_1 _0740_ (.A(net306),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[9] ),
    .X(_0189_));
 sg13g2_nand2_1 _0741_ (.Y(_0190_),
    .A(_0188_),
    .B(_0189_));
 sg13g2_nand3_1 _0742_ (.B(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ),
    .C(net113),
    .A(net383),
    .Y(_0191_));
 sg13g2_or2_1 _0743_ (.X(_0192_),
    .B(net384),
    .A(_0190_));
 sg13g2_inv_1 _0744_ (.Y(_0094_),
    .A(net385));
 sg13g2_nor2_2 _0745_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[1] ),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ),
    .Y(_0193_));
 sg13g2_nor2_1 _0746_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Done ),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_a22oi_1 _0747_ (.Y(_0015_),
    .B1(_0194_),
    .B2(_0192_),
    .A2(_0193_),
    .A1(_0128_));
 sg13g2_nand2_1 _0748_ (.Y(_0195_),
    .A(\TRNG_inst.U3_Main_controller.state[0] ),
    .B(net393));
 sg13g2_or2_1 _0749_ (.X(_0196_),
    .B(_0195_),
    .A(net114));
 sg13g2_nor2b_1 _0750_ (.A(\TRNG_inst.U3_Main_controller.state[0] ),
    .B_N(net360),
    .Y(_0197_));
 sg13g2_nand2_1 _0751_ (.Y(_0198_),
    .A(_0130_),
    .B(net360));
 sg13g2_nor2_1 _0752_ (.A(net114),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_o21ai_1 _0753_ (.B1(_0196_),
    .Y(_0016_),
    .A1(_0181_),
    .A2(_0199_));
 sg13g2_nor2_1 _0754_ (.A(_0129_),
    .B(net391),
    .Y(_0200_));
 sg13g2_a21oi_1 _0755_ (.A1(\TRNG_inst.U3_Main_controller.state[1] ),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0199_));
 sg13g2_o21ai_1 _0756_ (.B1(_0201_),
    .Y(_0202_),
    .A1(net335),
    .A2(_0130_));
 sg13g2_a21oi_1 _0757_ (.A1(_0182_),
    .A2(net361),
    .Y(_0017_),
    .B1(_0202_));
 sg13g2_and3_1 _0758_ (.X(_0203_),
    .A(_0127_),
    .B(\TRNG_inst.U3_Main_controller.cnt_bytes[1] ),
    .C(_0010_));
 sg13g2_nand2_1 _0759_ (.Y(_0204_),
    .A(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ),
    .B(net364));
 sg13g2_nor2_1 _0760_ (.A(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_nor2_2 _0761_ (.A(net110),
    .B(net109),
    .Y(_0206_));
 sg13g2_nor2b_1 _0762_ (.A(net114),
    .B_N(net335),
    .Y(_0207_));
 sg13g2_nand2b_1 _0763_ (.Y(_0208_),
    .B(\TRNG_inst.U3_Main_controller.state[2] ),
    .A_N(net114));
 sg13g2_nand2_1 _0764_ (.Y(_0209_),
    .A(\TRNG_inst.U3_Main_controller.state[0] ),
    .B(_0207_));
 sg13g2_a21oi_1 _0765_ (.A1(net242),
    .A2(net110),
    .Y(_0210_),
    .B1(net108));
 sg13g2_a22oi_1 _0766_ (.Y(_0211_),
    .B1(_0206_),
    .B2(\TRNG_inst.U3_Main_controller.tmp_reg[8] ),
    .A2(net109),
    .A1(\TRNG_inst.U3_Main_controller.tmp_reg[24] ));
 sg13g2_nor2_1 _0767_ (.A(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ),
    .B(net108),
    .Y(_0212_));
 sg13g2_a21oi_1 _0768_ (.A1(\TRNG_inst.U3_Main_controller.cnt_bytes[1] ),
    .A2(_0010_),
    .Y(_0213_),
    .B1(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ));
 sg13g2_o21ai_1 _0769_ (.B1(_0207_),
    .Y(_0214_),
    .A1(_0130_),
    .A2(_0010_));
 sg13g2_a21o_1 _0770_ (.A2(_0213_),
    .A1(_0212_),
    .B1(_0214_),
    .X(_0215_));
 sg13g2_a221oi_1 _0771_ (.B2(_0211_),
    .C1(net98),
    .B1(_0210_),
    .A1(_0152_),
    .Y(_0216_),
    .A2(net107));
 sg13g2_a21o_1 _0772_ (.A2(net98),
    .A1(net243),
    .B1(_0216_),
    .X(_0018_));
 sg13g2_a21oi_1 _0773_ (.A1(\TRNG_inst.U3_Main_controller.tmp_reg[17] ),
    .A2(net110),
    .Y(_0217_),
    .B1(net107));
 sg13g2_a22oi_1 _0774_ (.Y(_0218_),
    .B1(_0206_),
    .B2(net224),
    .A2(net109),
    .A1(\TRNG_inst.U3_Main_controller.tmp_reg[25] ));
 sg13g2_a221oi_1 _0775_ (.B2(_0218_),
    .C1(net99),
    .B1(_0217_),
    .A1(_0156_),
    .Y(_0219_),
    .A2(net107));
 sg13g2_a21o_1 _0776_ (.A2(net98),
    .A1(net232),
    .B1(_0219_),
    .X(_0019_));
 sg13g2_a21oi_1 _0777_ (.A1(\TRNG_inst.U3_Main_controller.tmp_reg[26] ),
    .A2(_0205_),
    .Y(_0220_),
    .B1(net108));
 sg13g2_a22oi_1 _0778_ (.Y(_0221_),
    .B1(_0206_),
    .B2(net263),
    .A2(net110),
    .A1(net254));
 sg13g2_a221oi_1 _0779_ (.B2(_0221_),
    .C1(_0215_),
    .B1(_0220_),
    .A1(_0160_),
    .Y(_0222_),
    .A2(net107));
 sg13g2_a21o_1 _0780_ (.A2(net98),
    .A1(net276),
    .B1(_0222_),
    .X(_0020_));
 sg13g2_a21oi_1 _0781_ (.A1(\TRNG_inst.U3_Main_controller.tmp_reg[27] ),
    .A2(net109),
    .Y(_0223_),
    .B1(net108));
 sg13g2_a22oi_1 _0782_ (.Y(_0224_),
    .B1(_0206_),
    .B2(\TRNG_inst.U3_Main_controller.tmp_reg[11] ),
    .A2(net110),
    .A1(\TRNG_inst.U3_Main_controller.tmp_reg[19] ));
 sg13g2_a221oi_1 _0783_ (.B2(_0224_),
    .C1(net99),
    .B1(_0223_),
    .A1(_0164_),
    .Y(_0225_),
    .A2(net107));
 sg13g2_a21o_1 _0784_ (.A2(net98),
    .A1(net285),
    .B1(_0225_),
    .X(_0021_));
 sg13g2_a21oi_1 _0785_ (.A1(\TRNG_inst.U3_Main_controller.tmp_reg[20] ),
    .A2(net110),
    .Y(_0226_),
    .B1(net106));
 sg13g2_a22oi_1 _0786_ (.Y(_0227_),
    .B1(_0206_),
    .B2(\TRNG_inst.U3_Main_controller.tmp_reg[12] ),
    .A2(net109),
    .A1(net234));
 sg13g2_a221oi_1 _0787_ (.B2(_0227_),
    .C1(net99),
    .B1(_0226_),
    .A1(_0168_),
    .Y(_0228_),
    .A2(net106));
 sg13g2_a21o_1 _0788_ (.A2(net98),
    .A1(net237),
    .B1(_0228_),
    .X(_0022_));
 sg13g2_a21oi_1 _0789_ (.A1(net259),
    .A2(_0203_),
    .Y(_0229_),
    .B1(net107));
 sg13g2_a22oi_1 _0790_ (.Y(_0230_),
    .B1(_0206_),
    .B2(net274),
    .A2(net109),
    .A1(net228));
 sg13g2_a221oi_1 _0791_ (.B2(_0230_),
    .C1(net99),
    .B1(_0229_),
    .A1(_0172_),
    .Y(_0231_),
    .A2(net107));
 sg13g2_a21o_1 _0792_ (.A2(net99),
    .A1(net288),
    .B1(_0231_),
    .X(_0023_));
 sg13g2_a21oi_1 _0793_ (.A1(net246),
    .A2(net110),
    .Y(_0232_),
    .B1(net106));
 sg13g2_a22oi_1 _0794_ (.Y(_0233_),
    .B1(_0206_),
    .B2(\TRNG_inst.U3_Main_controller.tmp_reg[14] ),
    .A2(net109),
    .A1(\TRNG_inst.U3_Main_controller.tmp_reg[30] ));
 sg13g2_a221oi_1 _0795_ (.B2(_0233_),
    .C1(net99),
    .B1(_0232_),
    .A1(_0176_),
    .Y(_0234_),
    .A2(net106));
 sg13g2_a21o_1 _0796_ (.A2(net98),
    .A1(net247),
    .B1(_0234_),
    .X(_0024_));
 sg13g2_a21oi_1 _0797_ (.A1(net230),
    .A2(net110),
    .Y(_0235_),
    .B1(net106));
 sg13g2_a22oi_1 _0798_ (.Y(_0236_),
    .B1(_0206_),
    .B2(\TRNG_inst.U3_Main_controller.tmp_reg[15] ),
    .A2(net109),
    .A1(\TRNG_inst.U3_Main_controller.tmp_reg[31] ));
 sg13g2_a221oi_1 _0799_ (.B2(_0236_),
    .C1(net99),
    .B1(_0235_),
    .A1(_0180_),
    .Y(_0237_),
    .A2(net107));
 sg13g2_a21o_1 _0800_ (.A2(net98),
    .A1(net209),
    .B1(net231),
    .X(_0025_));
 sg13g2_nand2_1 _0801_ (.Y(_0238_),
    .A(net112),
    .B(_0193_));
 sg13g2_nand3_1 _0802_ (.B(net204),
    .C(_0193_),
    .A(net113),
    .Y(_0239_));
 sg13g2_mux2_1 _0803_ (.A0(net243),
    .A1(net261),
    .S(_0239_),
    .X(_0026_));
 sg13g2_mux2_1 _0804_ (.A0(net232),
    .A1(net264),
    .S(net105),
    .X(_0027_));
 sg13g2_mux2_1 _0805_ (.A0(net276),
    .A1(net289),
    .S(net105),
    .X(_0028_));
 sg13g2_mux2_1 _0806_ (.A0(net285),
    .A1(net305),
    .S(net105),
    .X(_0029_));
 sg13g2_mux2_1 _0807_ (.A0(net237),
    .A1(net284),
    .S(net105),
    .X(_0030_));
 sg13g2_mux2_1 _0808_ (.A0(net288),
    .A1(net304),
    .S(net105),
    .X(_0031_));
 sg13g2_mux2_1 _0809_ (.A0(net247),
    .A1(net295),
    .S(net105),
    .X(_0032_));
 sg13g2_mux2_1 _0810_ (.A0(net209),
    .A1(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[7] ),
    .S(net105),
    .X(_0033_));
 sg13g2_nor3_1 _0811_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[3] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ),
    .Y(_0240_));
 sg13g2_nand2_1 _0812_ (.Y(_0241_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[4] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ));
 sg13g2_o21ai_1 _0813_ (.B1(_0137_),
    .Y(_0242_),
    .A1(_0240_),
    .A2(_0241_));
 sg13g2_and2_1 _0814_ (.A(net333),
    .B(net302),
    .X(_0243_));
 sg13g2_a21oi_2 _0815_ (.B1(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ),
    .Y(_0244_),
    .A2(_0243_),
    .A1(_0242_));
 sg13g2_a21o_2 _0816_ (.A2(_0243_),
    .A1(_0242_),
    .B1(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ),
    .X(_0245_));
 sg13g2_nand2_2 _0817_ (.Y(_0246_),
    .A(net349),
    .B(_0003_));
 sg13g2_nor2_1 _0818_ (.A(net372),
    .B(net350),
    .Y(_0247_));
 sg13g2_nand2b_2 _0819_ (.Y(_0248_),
    .B(_0134_),
    .A_N(_0246_));
 sg13g2_nor2_2 _0820_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ),
    .Y(_0249_));
 sg13g2_nand4_1 _0821_ (.B(_0245_),
    .C(_0247_),
    .A(_0008_),
    .Y(_0250_),
    .D(_0249_));
 sg13g2_nand2_1 _0822_ (.Y(_0251_),
    .A(net211),
    .B(_0250_));
 sg13g2_o21ai_1 _0823_ (.B1(net212),
    .Y(_0034_),
    .A1(_0140_),
    .A2(_0250_));
 sg13g2_xor2_1 _0824_ (.B(_0249_),
    .A(_0008_),
    .X(_0252_));
 sg13g2_nand3_1 _0825_ (.B(_0247_),
    .C(_0252_),
    .A(_0245_),
    .Y(_0253_));
 sg13g2_nand2_1 _0826_ (.Y(_0254_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ));
 sg13g2_nand2b_1 _0827_ (.Y(_0255_),
    .B(_0254_),
    .A_N(_0249_));
 sg13g2_or2_1 _0828_ (.X(_0256_),
    .B(_0255_),
    .A(net195));
 sg13g2_o21ai_1 _0829_ (.B1(net265),
    .Y(_0257_),
    .A1(_0253_),
    .A2(_0256_));
 sg13g2_nand3b_1 _0830_ (.B(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ),
    .Y(_0258_),
    .A_N(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ));
 sg13g2_o21ai_1 _0831_ (.B1(_0257_),
    .Y(_0035_),
    .A1(_0253_),
    .A2(_0258_));
 sg13g2_nand2_1 _0832_ (.Y(_0259_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .B(_0145_));
 sg13g2_o21ai_1 _0833_ (.B1(net225),
    .Y(_0260_),
    .A1(_0253_),
    .A2(_0259_));
 sg13g2_nor2_1 _0834_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ),
    .B(_0009_),
    .Y(_0261_));
 sg13g2_nand2_1 _0835_ (.Y(_0262_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .B(_0261_));
 sg13g2_o21ai_1 _0836_ (.B1(net226),
    .Y(_0036_),
    .A1(_0253_),
    .A2(_0262_));
 sg13g2_a21oi_1 _0837_ (.A1(_0008_),
    .A2(_0249_),
    .Y(_0263_),
    .B1(net195));
 sg13g2_nand2_1 _0838_ (.Y(_0264_),
    .A(_0255_),
    .B(_0263_));
 sg13g2_o21ai_1 _0839_ (.B1(net299),
    .Y(_0265_),
    .A1(_0253_),
    .A2(_0264_));
 sg13g2_nand3_1 _0840_ (.B(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ),
    .Y(_0266_));
 sg13g2_o21ai_1 _0841_ (.B1(_0265_),
    .Y(_0037_),
    .A1(_0253_),
    .A2(_0266_));
 sg13g2_o21ai_1 _0842_ (.B1(net239),
    .Y(_0267_),
    .A1(_0008_),
    .A2(_0253_));
 sg13g2_nand2b_1 _0843_ (.Y(_0268_),
    .B(_0261_),
    .A_N(_0253_));
 sg13g2_o21ai_1 _0844_ (.B1(net240),
    .Y(_0038_),
    .A1(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .A2(_0268_));
 sg13g2_or3_2 _0845_ (.A(_0244_),
    .B(_0248_),
    .C(_0252_),
    .X(_0269_));
 sg13g2_o21ai_1 _0846_ (.B1(net219),
    .Y(_0270_),
    .A1(_0256_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0847_ (.B1(_0270_),
    .Y(_0039_),
    .A1(_0258_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0848_ (.B1(net292),
    .Y(_0271_),
    .A1(_0259_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0849_ (.B1(net293),
    .Y(_0040_),
    .A1(_0262_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0850_ (.B1(net255),
    .Y(_0272_),
    .A1(_0264_),
    .A2(_0269_));
 sg13g2_o21ai_1 _0851_ (.B1(_0272_),
    .Y(_0041_),
    .A1(_0266_),
    .A2(_0269_));
 sg13g2_nor2_1 _0852_ (.A(net349),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ),
    .Y(_0273_));
 sg13g2_nand2_1 _0853_ (.Y(_0274_),
    .A(_0003_),
    .B(_0273_));
 sg13g2_o21ai_1 _0854_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0244_),
    .A2(_0248_));
 sg13g2_nor2_1 _0855_ (.A(_0008_),
    .B(_0254_),
    .Y(_0276_));
 sg13g2_nor2_1 _0856_ (.A(_0248_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nand3_1 _0857_ (.B(_0275_),
    .C(_0277_),
    .A(net195),
    .Y(_0278_));
 sg13g2_o21ai_1 _0858_ (.B1(_0278_),
    .Y(_0042_),
    .A1(_0145_),
    .A2(_0275_));
 sg13g2_nor2_1 _0859_ (.A(_0248_),
    .B(_0255_),
    .Y(_0279_));
 sg13g2_mux2_1 _0860_ (.A0(net380),
    .A1(_0279_),
    .S(_0275_),
    .X(_0043_));
 sg13g2_nand2b_1 _0861_ (.Y(_0280_),
    .B(_0275_),
    .A_N(_0254_));
 sg13g2_o21ai_1 _0862_ (.B1(_0277_),
    .Y(_0281_),
    .A1(_0144_),
    .A2(_0254_));
 sg13g2_a22oi_1 _0863_ (.Y(_0044_),
    .B1(_0281_),
    .B2(_0275_),
    .A2(_0280_),
    .A1(_0144_));
 sg13g2_and3_2 _0864_ (.X(_0282_),
    .A(net114),
    .B(\TRNG_inst.U3_Main_controller.state[0] ),
    .C(net360));
 sg13g2_nand3_1 _0865_ (.B(\TRNG_inst.U3_Main_controller.state[0] ),
    .C(_0001_),
    .A(net114),
    .Y(_0283_));
 sg13g2_nand4_1 _0866_ (.B(net222),
    .C(net308),
    .A(\TRNG_inst.U3_Main_controller.cnt_delay[6] ),
    .Y(_0284_),
    .D(net271));
 sg13g2_nand3_1 _0867_ (.B(\TRNG_inst.U3_Main_controller.cnt_delay[0] ),
    .C(\TRNG_inst.U3_Main_controller.cnt_delay[10] ),
    .A(\TRNG_inst.U3_Main_controller.cnt_delay[1] ),
    .Y(_0285_));
 sg13g2_nand4_1 _0868_ (.B(\TRNG_inst.U3_Main_controller.cnt_delay[8] ),
    .C(\TRNG_inst.U3_Main_controller.cnt_delay[3] ),
    .A(\TRNG_inst.U3_Main_controller.cnt_delay[9] ),
    .Y(_0286_),
    .D(\TRNG_inst.U3_Main_controller.cnt_delay[2] ));
 sg13g2_nor3_1 _0869_ (.A(_0284_),
    .B(_0285_),
    .C(_0286_),
    .Y(_0287_));
 sg13g2_nand2b_1 _0870_ (.Y(_0288_),
    .B(_0282_),
    .A_N(_0287_));
 sg13g2_inv_1 _0871_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_nor2_1 _0872_ (.A(_0195_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_and2_1 _0873_ (.A(_0282_),
    .B(_0287_),
    .X(_0291_));
 sg13g2_nand2_1 _0874_ (.Y(_0292_),
    .A(\TRNG_inst.U1_TRNG.o_data[0] ),
    .B(net103));
 sg13g2_o21ai_1 _0875_ (.B1(_0292_),
    .Y(_0045_),
    .A1(_0152_),
    .A2(net96));
 sg13g2_nand2_1 _0876_ (.Y(_0293_),
    .A(net206),
    .B(net103));
 sg13g2_o21ai_1 _0877_ (.B1(_0293_),
    .Y(_0046_),
    .A1(_0156_),
    .A2(net96));
 sg13g2_nand2_1 _0878_ (.Y(_0294_),
    .A(\TRNG_inst.U1_TRNG.o_data[2] ),
    .B(net103));
 sg13g2_o21ai_1 _0879_ (.B1(_0294_),
    .Y(_0047_),
    .A1(_0160_),
    .A2(net96));
 sg13g2_nand2_1 _0880_ (.Y(_0295_),
    .A(net198),
    .B(net103));
 sg13g2_o21ai_1 _0881_ (.B1(_0295_),
    .Y(_0048_),
    .A1(_0164_),
    .A2(net96));
 sg13g2_nand2_1 _0882_ (.Y(_0296_),
    .A(\TRNG_inst.U1_TRNG.o_data[4] ),
    .B(net103));
 sg13g2_o21ai_1 _0883_ (.B1(_0296_),
    .Y(_0049_),
    .A1(_0168_),
    .A2(net96));
 sg13g2_nand2_1 _0884_ (.Y(_0297_),
    .A(\TRNG_inst.U1_TRNG.o_data[5] ),
    .B(net103));
 sg13g2_o21ai_1 _0885_ (.B1(_0297_),
    .Y(_0050_),
    .A1(_0172_),
    .A2(net96));
 sg13g2_nand2_1 _0886_ (.Y(_0298_),
    .A(\TRNG_inst.U1_TRNG.o_data[6] ),
    .B(net103));
 sg13g2_o21ai_1 _0887_ (.B1(_0298_),
    .Y(_0051_),
    .A1(_0176_),
    .A2(net96));
 sg13g2_nand2_1 _0888_ (.Y(_0299_),
    .A(net194),
    .B(net100));
 sg13g2_o21ai_1 _0889_ (.B1(_0299_),
    .Y(_0052_),
    .A1(_0180_),
    .A2(net93));
 sg13g2_nand2_1 _0890_ (.Y(_0300_),
    .A(\TRNG_inst.U1_TRNG.o_data[8] ),
    .B(net101));
 sg13g2_o21ai_1 _0891_ (.B1(_0300_),
    .Y(_0053_),
    .A1(_0151_),
    .A2(net94));
 sg13g2_nand2_1 _0892_ (.Y(_0301_),
    .A(net197),
    .B(net101));
 sg13g2_o21ai_1 _0893_ (.B1(_0301_),
    .Y(_0054_),
    .A1(_0155_),
    .A2(net94));
 sg13g2_nand2_1 _0894_ (.Y(_0302_),
    .A(\TRNG_inst.U1_TRNG.o_data[10] ),
    .B(net100));
 sg13g2_o21ai_1 _0895_ (.B1(_0302_),
    .Y(_0055_),
    .A1(_0159_),
    .A2(net93));
 sg13g2_nand2_1 _0896_ (.Y(_0303_),
    .A(\TRNG_inst.U1_TRNG.o_data[11] ),
    .B(net100));
 sg13g2_o21ai_1 _0897_ (.B1(_0303_),
    .Y(_0056_),
    .A1(_0163_),
    .A2(net93));
 sg13g2_nand2_1 _0898_ (.Y(_0304_),
    .A(\TRNG_inst.U1_TRNG.o_data[12] ),
    .B(net100));
 sg13g2_o21ai_1 _0899_ (.B1(_0304_),
    .Y(_0057_),
    .A1(_0167_),
    .A2(net93));
 sg13g2_nand2_1 _0900_ (.Y(_0305_),
    .A(\TRNG_inst.U1_TRNG.o_data[13] ),
    .B(net101));
 sg13g2_o21ai_1 _0901_ (.B1(_0305_),
    .Y(_0058_),
    .A1(_0171_),
    .A2(net94));
 sg13g2_nand2_1 _0902_ (.Y(_0306_),
    .A(\TRNG_inst.U1_TRNG.o_data[14] ),
    .B(net101));
 sg13g2_o21ai_1 _0903_ (.B1(_0306_),
    .Y(_0059_),
    .A1(_0175_),
    .A2(net94));
 sg13g2_nand2_1 _0904_ (.Y(_0307_),
    .A(net201),
    .B(net101));
 sg13g2_o21ai_1 _0905_ (.B1(_0307_),
    .Y(_0060_),
    .A1(_0179_),
    .A2(net94));
 sg13g2_nand2_1 _0906_ (.Y(_0308_),
    .A(\TRNG_inst.U1_TRNG.o_data[16] ),
    .B(net102));
 sg13g2_o21ai_1 _0907_ (.B1(_0308_),
    .Y(_0061_),
    .A1(_0150_),
    .A2(net97));
 sg13g2_nand2_1 _0908_ (.Y(_0309_),
    .A(\TRNG_inst.U1_TRNG.o_data[17] ),
    .B(net102));
 sg13g2_o21ai_1 _0909_ (.B1(_0309_),
    .Y(_0062_),
    .A1(_0154_),
    .A2(net95));
 sg13g2_nand2_1 _0910_ (.Y(_0310_),
    .A(net235),
    .B(net100));
 sg13g2_o21ai_1 _0911_ (.B1(_0310_),
    .Y(_0063_),
    .A1(_0158_),
    .A2(net93));
 sg13g2_nand2_1 _0912_ (.Y(_0311_),
    .A(\TRNG_inst.U1_TRNG.o_data[19] ),
    .B(net100));
 sg13g2_o21ai_1 _0913_ (.B1(_0311_),
    .Y(_0064_),
    .A1(_0162_),
    .A2(net93));
 sg13g2_nand2_1 _0914_ (.Y(_0312_),
    .A(\TRNG_inst.U1_TRNG.o_data[20] ),
    .B(net100));
 sg13g2_o21ai_1 _0915_ (.B1(_0312_),
    .Y(_0065_),
    .A1(_0166_),
    .A2(net93));
 sg13g2_nand2_1 _0916_ (.Y(_0313_),
    .A(\TRNG_inst.U1_TRNG.o_data[21] ),
    .B(net102));
 sg13g2_o21ai_1 _0917_ (.B1(_0313_),
    .Y(_0066_),
    .A1(_0170_),
    .A2(net95));
 sg13g2_nand2_1 _0918_ (.Y(_0314_),
    .A(\TRNG_inst.U1_TRNG.o_data[22] ),
    .B(net102));
 sg13g2_o21ai_1 _0919_ (.B1(_0314_),
    .Y(_0067_),
    .A1(_0174_),
    .A2(net95));
 sg13g2_nand2_1 _0920_ (.Y(_0315_),
    .A(\TRNG_inst.U1_TRNG.o_data[23] ),
    .B(net100));
 sg13g2_o21ai_1 _0921_ (.B1(_0315_),
    .Y(_0068_),
    .A1(_0178_),
    .A2(net93));
 sg13g2_nand2_1 _0922_ (.Y(_0316_),
    .A(net217),
    .B(net101));
 sg13g2_o21ai_1 _0923_ (.B1(_0316_),
    .Y(_0069_),
    .A1(_0149_),
    .A2(net94));
 sg13g2_nand2_1 _0924_ (.Y(_0317_),
    .A(\TRNG_inst.U1_TRNG.o_data[25] ),
    .B(net101));
 sg13g2_o21ai_1 _0925_ (.B1(_0317_),
    .Y(_0070_),
    .A1(_0153_),
    .A2(net94));
 sg13g2_nand2_1 _0926_ (.Y(_0318_),
    .A(net215),
    .B(net104));
 sg13g2_o21ai_1 _0927_ (.B1(_0318_),
    .Y(_0071_),
    .A1(_0157_),
    .A2(net97));
 sg13g2_nand2_1 _0928_ (.Y(_0319_),
    .A(\TRNG_inst.U1_TRNG.o_data[27] ),
    .B(net104));
 sg13g2_o21ai_1 _0929_ (.B1(_0319_),
    .Y(_0072_),
    .A1(_0161_),
    .A2(net97));
 sg13g2_nand2_1 _0930_ (.Y(_0320_),
    .A(\TRNG_inst.U1_TRNG.o_data[28] ),
    .B(net104));
 sg13g2_o21ai_1 _0931_ (.B1(_0320_),
    .Y(_0073_),
    .A1(_0165_),
    .A2(net95));
 sg13g2_nand2_1 _0932_ (.Y(_0321_),
    .A(net199),
    .B(net103));
 sg13g2_o21ai_1 _0933_ (.B1(_0321_),
    .Y(_0074_),
    .A1(_0169_),
    .A2(net96));
 sg13g2_nand2_1 _0934_ (.Y(_0322_),
    .A(\TRNG_inst.U1_TRNG.o_data[30] ),
    .B(net102));
 sg13g2_o21ai_1 _0935_ (.B1(_0322_),
    .Y(_0075_),
    .A1(_0173_),
    .A2(net95));
 sg13g2_nand2_1 _0936_ (.Y(_0323_),
    .A(\TRNG_inst.U1_TRNG.o_data[31] ),
    .B(net101));
 sg13g2_o21ai_1 _0937_ (.B1(_0323_),
    .Y(_0076_),
    .A1(_0177_),
    .A2(net94));
 sg13g2_nand3b_1 _0938_ (.B(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ),
    .C(net112),
    .Y(_0324_),
    .A_N(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[1] ));
 sg13g2_a21oi_1 _0939_ (.A1(_0147_),
    .A2(_0324_),
    .Y(_0077_),
    .B1(_0193_));
 sg13g2_nand2_1 _0940_ (.Y(_0325_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ),
    .B(_0003_));
 sg13g2_nor3_1 _0941_ (.A(_0134_),
    .B(_0244_),
    .C(net350),
    .Y(_0107_));
 sg13g2_o21ai_1 _0942_ (.B1(_0273_),
    .Y(_0326_),
    .A1(net357),
    .A2(net111));
 sg13g2_o21ai_1 _0943_ (.B1(net358),
    .Y(_0327_),
    .A1(\TRNG_inst.U2_UART_interface.RX_part.r_RX_DV ),
    .A2(net351));
 sg13g2_inv_1 _0944_ (.Y(_0078_),
    .A(net359));
 sg13g2_a22oi_1 _0945_ (.Y(_0328_),
    .B1(_0289_),
    .B2(net189),
    .A2(_0283_),
    .A1(\TRNG_inst.U3_Main_controller.cnt_delay[0] ));
 sg13g2_inv_1 _0946_ (.Y(_0079_),
    .A(net190));
 sg13g2_nand3_1 _0947_ (.B(\TRNG_inst.U3_Main_controller.cnt_delay[0] ),
    .C(_0282_),
    .A(net376),
    .Y(_0329_));
 sg13g2_a21o_1 _0948_ (.A2(_0282_),
    .A1(\TRNG_inst.U3_Main_controller.cnt_delay[0] ),
    .B1(net376),
    .X(_0330_));
 sg13g2_and2_1 _0949_ (.A(_0329_),
    .B(net377),
    .X(_0080_));
 sg13g2_and4_1 _0950_ (.A(net250),
    .B(\TRNG_inst.U3_Main_controller.cnt_delay[1] ),
    .C(\TRNG_inst.U3_Main_controller.cnt_delay[0] ),
    .D(_0282_),
    .X(_0331_));
 sg13g2_xnor2_1 _0951_ (.Y(_0081_),
    .A(net250),
    .B(_0329_));
 sg13g2_nand2_1 _0952_ (.Y(_0332_),
    .A(net311),
    .B(_0331_));
 sg13g2_xor2_1 _0953_ (.B(_0331_),
    .A(net311),
    .X(_0082_));
 sg13g2_and3_1 _0954_ (.X(_0333_),
    .A(net271),
    .B(\TRNG_inst.U3_Main_controller.cnt_delay[3] ),
    .C(_0331_));
 sg13g2_xnor2_1 _0955_ (.Y(_0083_),
    .A(net271),
    .B(_0332_));
 sg13g2_xor2_1 _0956_ (.B(_0333_),
    .A(net308),
    .X(_0084_));
 sg13g2_nand3_1 _0957_ (.B(net308),
    .C(_0333_),
    .A(net375),
    .Y(_0334_));
 sg13g2_a21o_1 _0958_ (.A2(_0333_),
    .A1(net308),
    .B1(net375),
    .X(_0335_));
 sg13g2_and2_1 _0959_ (.A(_0334_),
    .B(_0335_),
    .X(_0085_));
 sg13g2_nor2_2 _0960_ (.A(_0284_),
    .B(_0332_),
    .Y(_0336_));
 sg13g2_a21oi_1 _0961_ (.A1(_0146_),
    .A2(_0334_),
    .Y(_0086_),
    .B1(_0336_));
 sg13g2_xor2_1 _0962_ (.B(_0336_),
    .A(net316),
    .X(_0087_));
 sg13g2_nand3_1 _0963_ (.B(net316),
    .C(_0336_),
    .A(net374),
    .Y(_0337_));
 sg13g2_a21o_1 _0964_ (.A2(_0336_),
    .A1(net316),
    .B1(net374),
    .X(_0338_));
 sg13g2_and2_1 _0965_ (.A(_0337_),
    .B(_0338_),
    .X(_0088_));
 sg13g2_xnor2_1 _0966_ (.Y(_0089_),
    .A(net257),
    .B(_0337_));
 sg13g2_nor3_1 _0967_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[1] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[3] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[2] ),
    .Y(_0339_));
 sg13g2_nand4_1 _0968_ (.B(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[0] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[4] ),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_DV ),
    .Y(_0340_),
    .D(_0339_));
 sg13g2_nor4_2 _0969_ (.A(_0148_),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[7] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[6] ),
    .Y(_0341_),
    .D(_0340_));
 sg13g2_o21ai_1 _0970_ (.B1(_0288_),
    .Y(_0342_),
    .A1(_0196_),
    .A2(_0341_));
 sg13g2_or2_1 _0971_ (.X(_0343_),
    .B(_0342_),
    .A(_0212_));
 sg13g2_nor3_1 _0972_ (.A(_0207_),
    .B(_0282_),
    .C(_0342_),
    .Y(_0344_));
 sg13g2_a21oi_1 _0973_ (.A1(_0129_),
    .A2(_0343_),
    .Y(_0090_),
    .B1(_0344_));
 sg13g2_nand2_1 _0974_ (.Y(_0345_),
    .A(_0196_),
    .B(net106));
 sg13g2_a21oi_1 _0975_ (.A1(net114),
    .A2(_0197_),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_o21ai_1 _0976_ (.B1(_0288_),
    .Y(_0091_),
    .A1(_0343_),
    .A2(net388));
 sg13g2_nor2_1 _0977_ (.A(net114),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_RX_DV ),
    .Y(_0347_));
 sg13g2_nor2_1 _0978_ (.A(_0198_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_or3_1 _0979_ (.A(_0200_),
    .B(_0343_),
    .C(_0348_),
    .X(_0092_));
 sg13g2_mux2_1 _0980_ (.A0(net261),
    .A1(net264),
    .S(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .X(_0349_));
 sg13g2_nand2_1 _0981_ (.Y(_0350_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .B(net338));
 sg13g2_inv_1 _0982_ (.Y(_0351_),
    .A(_0350_));
 sg13g2_nor2b_1 _0983_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .B_N(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[2] ),
    .Y(_0352_));
 sg13g2_a21oi_1 _0984_ (.A1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .A2(net305),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_a21oi_1 _0985_ (.A1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ),
    .A2(_0353_),
    .Y(_0354_),
    .B1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[2] ));
 sg13g2_o21ai_1 _0986_ (.B1(_0354_),
    .Y(_0355_),
    .A1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ),
    .A2(_0349_));
 sg13g2_mux4_1 _0987_ (.S0(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .A0(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[4] ),
    .A1(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[5] ),
    .A2(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[6] ),
    .A3(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[7] ),
    .S1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ),
    .X(_0356_));
 sg13g2_nand3b_1 _0988_ (.B(net112),
    .C(net383),
    .Y(_0357_),
    .A_N(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ));
 sg13g2_a21oi_1 _0989_ (.A1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[2] ),
    .A2(_0356_),
    .Y(_0358_),
    .B1(_0357_));
 sg13g2_o21ai_1 _0990_ (.B1(_0324_),
    .Y(_0359_),
    .A1(net112),
    .A2(net327));
 sg13g2_a21oi_1 _0991_ (.A1(_0355_),
    .A2(_0358_),
    .Y(_0093_),
    .B1(net328));
 sg13g2_a21oi_1 _0992_ (.A1(_0188_),
    .A2(_0189_),
    .Y(_0360_),
    .B1(_0191_));
 sg13g2_nand2b_1 _0993_ (.Y(_0361_),
    .B(_0190_),
    .A_N(net384));
 sg13g2_nor2_1 _0994_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .Y(_0362_));
 sg13g2_or2_1 _0995_ (.X(_0363_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ));
 sg13g2_nand2_1 _0996_ (.Y(_0364_),
    .A(net318),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ));
 sg13g2_nand4_1 _0997_ (.B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ),
    .C(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[8] ),
    .Y(_0365_),
    .D(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ));
 sg13g2_a21oi_1 _0998_ (.A1(_0362_),
    .A2(_0364_),
    .Y(_0366_),
    .B1(_0365_));
 sg13g2_nand2_1 _0999_ (.Y(_0367_),
    .A(net341),
    .B(net322));
 sg13g2_and3_1 _1000_ (.X(_0368_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[8] ),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ),
    .C(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ));
 sg13g2_nand2b_1 _1001_ (.Y(_0369_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[1] ),
    .A_N(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ));
 sg13g2_nor4_1 _1002_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ),
    .B(_0363_),
    .C(_0365_),
    .D(_0369_),
    .Y(_0370_));
 sg13g2_nor4_2 _1003_ (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[9] ),
    .B(_0366_),
    .C(_0368_),
    .Y(_0371_),
    .D(_0370_));
 sg13g2_o21ai_1 _1004_ (.B1(_0357_),
    .Y(_0372_),
    .A1(_0324_),
    .A2(_0371_));
 sg13g2_nand2b_1 _1005_ (.Y(_0095_),
    .B(_0361_),
    .A_N(_0372_));
 sg13g2_or4_1 _1006_ (.A(net381),
    .B(_0350_),
    .C(_0357_),
    .D(_0371_),
    .X(_0373_));
 sg13g2_nand2b_1 _1007_ (.Y(_0374_),
    .B(_0371_),
    .A_N(_0324_));
 sg13g2_nand4_1 _1008_ (.B(_0361_),
    .C(_0373_),
    .A(net105),
    .Y(_0096_),
    .D(_0374_));
 sg13g2_nand2b_1 _1009_ (.Y(_0375_),
    .B(net343),
    .A_N(net113));
 sg13g2_nor2b_1 _1010_ (.A(_0193_),
    .B_N(net112),
    .Y(_0376_));
 sg13g2_o21ai_1 _1011_ (.B1(_0376_),
    .Y(_0377_),
    .A1(_0360_),
    .A2(_0371_));
 sg13g2_and3_1 _1012_ (.X(_0378_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[1] ),
    .C(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ));
 sg13g2_nand2_1 _1013_ (.Y(_0379_),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .B(_0378_));
 sg13g2_nand4_1 _1014_ (.B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ),
    .C(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ),
    .Y(_0380_),
    .D(_0378_));
 sg13g2_nor3_1 _1015_ (.A(_0004_),
    .B(_0367_),
    .C(_0380_),
    .Y(_0381_));
 sg13g2_xnor2_1 _1016_ (.Y(_0382_),
    .A(net343),
    .B(_0381_));
 sg13g2_o21ai_1 _1017_ (.B1(_0375_),
    .Y(_0097_),
    .A1(net92),
    .A2(_0382_));
 sg13g2_nand2b_1 _1018_ (.Y(_0383_),
    .B(net306),
    .A_N(net112));
 sg13g2_o21ai_1 _1019_ (.B1(_0004_),
    .Y(_0384_),
    .A1(_0367_),
    .A2(_0380_));
 sg13g2_nand2b_1 _1020_ (.Y(_0385_),
    .B(_0384_),
    .A_N(_0381_));
 sg13g2_o21ai_1 _1021_ (.B1(_0383_),
    .Y(_0098_),
    .A1(net92),
    .A2(_0385_));
 sg13g2_nand2b_1 _1022_ (.Y(_0386_),
    .B(net322),
    .A_N(net112));
 sg13g2_nor2_1 _1023_ (.A(_0007_),
    .B(_0380_),
    .Y(_0387_));
 sg13g2_xor2_1 _1024_ (.B(_0387_),
    .A(_0005_),
    .X(_0388_));
 sg13g2_o21ai_1 _1025_ (.B1(_0386_),
    .Y(_0099_),
    .A1(net92),
    .A2(_0388_));
 sg13g2_nand2b_1 _1026_ (.Y(_0389_),
    .B(net341),
    .A_N(net324));
 sg13g2_xnor2_1 _1027_ (.Y(_0390_),
    .A(_0007_),
    .B(_0380_));
 sg13g2_o21ai_1 _1028_ (.B1(_0389_),
    .Y(_0100_),
    .A1(net92),
    .A2(_0390_));
 sg13g2_nand2b_1 _1029_ (.Y(_0391_),
    .B(net330),
    .A_N(net324));
 sg13g2_o21ai_1 _1030_ (.B1(_0141_),
    .Y(_0392_),
    .A1(_0142_),
    .A2(_0379_));
 sg13g2_nand2_1 _1031_ (.Y(_0393_),
    .A(_0380_),
    .B(_0392_));
 sg13g2_o21ai_1 _1032_ (.B1(_0391_),
    .Y(_0101_),
    .A1(net92),
    .A2(_0393_));
 sg13g2_nand2b_1 _1033_ (.Y(_0394_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ),
    .A_N(net324));
 sg13g2_xnor2_1 _1034_ (.Y(_0395_),
    .A(_0142_),
    .B(_0379_));
 sg13g2_o21ai_1 _1035_ (.B1(net325),
    .Y(_0102_),
    .A1(_0377_),
    .A2(_0395_));
 sg13g2_nand2b_1 _1036_ (.Y(_0396_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ),
    .A_N(net113));
 sg13g2_xor2_1 _1037_ (.B(_0378_),
    .A(net352),
    .X(_0397_));
 sg13g2_o21ai_1 _1038_ (.B1(_0396_),
    .Y(_0103_),
    .A1(net92),
    .A2(net353));
 sg13g2_nand2b_1 _1039_ (.Y(_0398_),
    .B(net355),
    .A_N(net113));
 sg13g2_xor2_1 _1040_ (.B(_0364_),
    .A(net355),
    .X(_0399_));
 sg13g2_o21ai_1 _1041_ (.B1(_0398_),
    .Y(_0104_),
    .A1(net92),
    .A2(_0399_));
 sg13g2_nand2b_1 _1042_ (.Y(_0400_),
    .B(net318),
    .A_N(net113));
 sg13g2_nand2_1 _1043_ (.Y(_0401_),
    .A(_0184_),
    .B(_0364_));
 sg13g2_o21ai_1 _1044_ (.B1(net319),
    .Y(_0105_),
    .A1(net92),
    .A2(_0401_));
 sg13g2_nand2b_1 _1045_ (.Y(_0402_),
    .B(net346),
    .A_N(net113));
 sg13g2_o21ai_1 _1046_ (.B1(_0402_),
    .Y(_0106_),
    .A1(net346),
    .A2(_0377_));
 sg13g2_nor2_2 _1047_ (.A(_0245_),
    .B(net350),
    .Y(_0403_));
 sg13g2_inv_1 _1048_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_nand3b_1 _1049_ (.B(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ),
    .C(net111),
    .Y(_0405_),
    .A_N(net349));
 sg13g2_inv_1 _1050_ (.Y(_0406_),
    .A(_0405_));
 sg13g2_nor4_2 _1051_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[8] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ),
    .Y(_0407_),
    .D(_0139_));
 sg13g2_nand2_1 _1052_ (.Y(_0408_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[4] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[3] ));
 sg13g2_nand2_1 _1053_ (.Y(_0409_),
    .A(net302),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[6] ));
 sg13g2_nor4_2 _1054_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ),
    .C(_0408_),
    .Y(_0410_),
    .D(_0409_));
 sg13g2_and2_1 _1055_ (.A(_0407_),
    .B(_0410_),
    .X(_0411_));
 sg13g2_nand3_1 _1056_ (.B(_0406_),
    .C(_0411_),
    .A(net336),
    .Y(_0412_));
 sg13g2_nand3_1 _1057_ (.B(_0404_),
    .C(_0412_),
    .A(_0248_),
    .Y(_0108_));
 sg13g2_nand3_1 _1058_ (.B(_0247_),
    .C(_0276_),
    .A(_0245_),
    .Y(_0413_));
 sg13g2_nor2_1 _1059_ (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ),
    .B(_0274_),
    .Y(_0414_));
 sg13g2_nor2_1 _1060_ (.A(_0405_),
    .B(_0411_),
    .Y(_0415_));
 sg13g2_nor2_1 _1061_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nand2_1 _1062_ (.Y(_0417_),
    .A(net372),
    .B(_0403_));
 sg13g2_nand3_1 _1063_ (.B(_0416_),
    .C(_0417_),
    .A(_0413_),
    .Y(_0109_));
 sg13g2_nor2_1 _1064_ (.A(_0140_),
    .B(_0405_),
    .Y(_0418_));
 sg13g2_and3_1 _1065_ (.X(_0419_),
    .A(_0407_),
    .B(_0410_),
    .C(_0418_));
 sg13g2_nand3_1 _1066_ (.B(_0410_),
    .C(_0418_),
    .A(_0407_),
    .Y(_0420_));
 sg13g2_nor2_2 _1067_ (.A(_0135_),
    .B(_0419_),
    .Y(_0421_));
 sg13g2_nand2_1 _1068_ (.Y(_0422_),
    .A(net111),
    .B(_0420_));
 sg13g2_and3_1 _1069_ (.X(_0423_),
    .A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ),
    .B(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ),
    .C(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[0] ));
 sg13g2_nand2b_2 _1070_ (.Y(_0424_),
    .B(_0423_),
    .A_N(_0408_));
 sg13g2_nor3_2 _1071_ (.A(_0135_),
    .B(_0419_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_nor3_2 _1072_ (.A(_0138_),
    .B(_0409_),
    .C(_0424_),
    .Y(_0426_));
 sg13g2_nand4_1 _1073_ (.B(net333),
    .C(_0420_),
    .A(net111),
    .Y(_0427_),
    .D(_0426_));
 sg13g2_xor2_1 _1074_ (.B(_0427_),
    .A(net370),
    .X(_0428_));
 sg13g2_a21oi_1 _1075_ (.A1(net111),
    .A2(_0405_),
    .Y(_0110_),
    .B1(_0428_));
 sg13g2_a21oi_1 _1076_ (.A1(_0421_),
    .A2(_0426_),
    .Y(_0429_),
    .B1(net333));
 sg13g2_a22oi_1 _1077_ (.Y(_0430_),
    .B1(_0405_),
    .B2(_0245_),
    .A2(_0325_),
    .A1(_0246_));
 sg13g2_nor2_1 _1078_ (.A(_0422_),
    .B(_0430_),
    .Y(_0431_));
 sg13g2_o21ai_1 _1079_ (.B1(_0427_),
    .Y(_0432_),
    .A1(_0422_),
    .A2(_0430_));
 sg13g2_nor2_1 _1080_ (.A(net334),
    .B(_0432_),
    .Y(_0111_));
 sg13g2_or4_1 _1081_ (.A(_0135_),
    .B(_0138_),
    .C(_0419_),
    .D(_0424_),
    .X(_0433_));
 sg13g2_or2_1 _1082_ (.X(_0434_),
    .B(_0433_),
    .A(_0137_));
 sg13g2_nor3_2 _1083_ (.A(_0403_),
    .B(_0415_),
    .C(_0422_),
    .Y(_0435_));
 sg13g2_a221oi_1 _1084_ (.B2(_0136_),
    .C1(_0435_),
    .B1(_0434_),
    .A1(_0421_),
    .Y(_0112_),
    .A2(_0426_));
 sg13g2_xnor2_1 _1085_ (.Y(_0436_),
    .A(_0137_),
    .B(_0433_));
 sg13g2_nor2_1 _1086_ (.A(_0435_),
    .B(_0436_),
    .Y(_0113_));
 sg13g2_xnor2_1 _1087_ (.Y(_0437_),
    .A(net363),
    .B(_0425_));
 sg13g2_nor2_1 _1088_ (.A(_0431_),
    .B(_0437_),
    .Y(_0114_));
 sg13g2_nor3_1 _1089_ (.A(_0135_),
    .B(_0139_),
    .C(_0419_),
    .Y(_0438_));
 sg13g2_nand4_1 _1090_ (.B(net366),
    .C(net345),
    .A(net111),
    .Y(_0439_),
    .D(_0420_));
 sg13g2_and4_1 _1091_ (.A(net111),
    .B(net280),
    .C(_0420_),
    .D(_0423_),
    .X(_0440_));
 sg13g2_nor2_1 _1092_ (.A(net321),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_nor3_1 _1093_ (.A(_0425_),
    .B(_0435_),
    .C(_0441_),
    .Y(_0115_));
 sg13g2_a21oi_1 _1094_ (.A1(_0421_),
    .A2(_0423_),
    .Y(_0442_),
    .B1(net280));
 sg13g2_nor3_1 _1095_ (.A(_0435_),
    .B(_0440_),
    .C(net281),
    .Y(_0116_));
 sg13g2_xor2_1 _1096_ (.B(_0439_),
    .A(net369),
    .X(_0443_));
 sg13g2_nor2_1 _1097_ (.A(_0431_),
    .B(_0443_),
    .Y(_0117_));
 sg13g2_xnor2_1 _1098_ (.Y(_0444_),
    .A(net366),
    .B(_0438_));
 sg13g2_nor2_1 _1099_ (.A(_0435_),
    .B(_0444_),
    .Y(_0118_));
 sg13g2_nor2_1 _1100_ (.A(net345),
    .B(_0421_),
    .Y(_0445_));
 sg13g2_nor3_1 _1101_ (.A(_0431_),
    .B(_0438_),
    .C(_0445_),
    .Y(_0119_));
 sg13g2_nor3_1 _1102_ (.A(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ),
    .B(\TRNG_inst.U3_Main_controller.cnt_bytes[1] ),
    .C(_0010_),
    .Y(_0446_));
 sg13g2_nand2b_1 _1103_ (.Y(_0447_),
    .B(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Done ),
    .A_N(net202));
 sg13g2_nor4_2 _1104_ (.A(net367),
    .B(net108),
    .C(_0446_),
    .Y(_0448_),
    .D(_0447_));
 sg13g2_a21oi_1 _1105_ (.A1(_0201_),
    .A2(net108),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_a21oi_1 _1106_ (.A1(_0143_),
    .A2(_0208_),
    .Y(_0120_),
    .B1(_0449_));
 sg13g2_o21ai_1 _1107_ (.B1(_0238_),
    .Y(_0450_),
    .A1(_0357_),
    .A2(_0371_));
 sg13g2_a21oi_1 _1108_ (.A1(_0133_),
    .A2(_0351_),
    .Y(_0451_),
    .B1(_0357_));
 sg13g2_nand3_1 _1109_ (.B(_0450_),
    .C(_0451_),
    .A(net191),
    .Y(_0452_));
 sg13g2_o21ai_1 _1110_ (.B1(net192),
    .Y(_0121_),
    .A1(_0132_),
    .A2(_0450_));
 sg13g2_nand2_1 _1111_ (.Y(_0453_),
    .A(_0351_),
    .B(_0450_));
 sg13g2_a21oi_1 _1112_ (.A1(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ),
    .A2(_0450_),
    .Y(_0454_),
    .B1(net338));
 sg13g2_a221oi_1 _1113_ (.B2(_0450_),
    .C1(net339),
    .B1(_0351_),
    .A1(net112),
    .Y(_0122_),
    .A2(_0193_));
 sg13g2_o21ai_1 _1114_ (.B1(_0451_),
    .Y(_0455_),
    .A1(_0131_),
    .A2(_0350_));
 sg13g2_a22oi_1 _1115_ (.Y(_0123_),
    .B1(_0455_),
    .B2(_0450_),
    .A2(_0453_),
    .A1(_0131_));
 sg13g2_nand2b_1 _1116_ (.Y(_0456_),
    .B(_0447_),
    .A_N(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ));
 sg13g2_nor2_1 _1117_ (.A(_0446_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _1118_ (.A(net106),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nand2_1 _1119_ (.Y(_0459_),
    .A(net186),
    .B(_0448_));
 sg13g2_o21ai_1 _1120_ (.B1(net187),
    .Y(_0124_),
    .A1(_0127_),
    .A2(_0458_));
 sg13g2_a21oi_1 _1121_ (.A1(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ),
    .A2(net364),
    .Y(_0460_),
    .B1(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ));
 sg13g2_o21ai_1 _1122_ (.B1(_0460_),
    .Y(_0461_),
    .A1(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ),
    .A2(net364));
 sg13g2_nor2_1 _1123_ (.A(net364),
    .B(_0458_),
    .Y(_0462_));
 sg13g2_a21oi_1 _1124_ (.A1(_0458_),
    .A2(_0461_),
    .Y(_0125_),
    .B1(_0462_));
 sg13g2_xor2_1 _1125_ (.B(_0204_),
    .A(_0010_),
    .X(_0463_));
 sg13g2_a22oi_1 _1126_ (.Y(_0464_),
    .B1(_0448_),
    .B2(_0463_),
    .A2(net106),
    .A1(net367));
 sg13g2_inv_1 _1127_ (.Y(_0126_),
    .A(net368));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net42),
    .D(net208),
    .Q_N(_0562_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Done ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net89),
    .D(net270),
    .Q_N(_0561_),
    .Q(\TRNG_inst.U3_Main_controller.led ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net88),
    .D(net362),
    .Q_N(_0560_),
    .Q(\TRNG_inst.U1_TRNG.i_rst ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net87),
    .D(net244),
    .Q_N(_0559_),
    .Q(\TRNG_inst.TX_Byte[0] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net86),
    .D(net233),
    .Q_N(_0558_),
    .Q(\TRNG_inst.TX_Byte[1] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net85),
    .D(net277),
    .Q_N(_0557_),
    .Q(\TRNG_inst.TX_Byte[2] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net84),
    .D(net286),
    .Q_N(_0556_),
    .Q(\TRNG_inst.TX_Byte[3] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net83),
    .D(net238),
    .Q_N(_0555_),
    .Q(\TRNG_inst.TX_Byte[4] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net82),
    .D(_0023_),
    .Q_N(_0554_),
    .Q(\TRNG_inst.TX_Byte[5] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net81),
    .D(net248),
    .Q_N(_0553_),
    .Q(\TRNG_inst.TX_Byte[6] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net80),
    .D(_0025_),
    .Q_N(_0552_),
    .Q(\TRNG_inst.TX_Byte[7] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net79),
    .D(_0026_),
    .Q_N(_0551_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[0] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net78),
    .D(_0027_),
    .Q_N(_0550_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[1] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net77),
    .D(_0028_),
    .Q_N(_0549_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[2] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net76),
    .D(_0029_),
    .Q_N(_0548_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[3] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net75),
    .D(_0030_),
    .Q_N(_0547_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[4] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net74),
    .D(_0031_),
    .Q_N(_0546_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[5] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net73),
    .D(_0032_),
    .Q_N(_0545_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[6] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net43),
    .D(net210),
    .Q_N(_0563_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[7] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net48),
    .D(net166),
    .Q_N(_0009_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net72),
    .D(net2),
    .Q_N(_0544_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data_R ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net71),
    .D(net213),
    .Q_N(_0543_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[0] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net70),
    .D(net266),
    .Q_N(_0542_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[1] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net69),
    .D(net227),
    .Q_N(_0541_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[2] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net68),
    .D(net300),
    .Q_N(_0540_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[3] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net67),
    .D(net241),
    .Q_N(_0539_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[4] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net66),
    .D(net220),
    .Q_N(_0538_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[5] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net65),
    .D(net294),
    .Q_N(_0537_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[6] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net64),
    .D(net256),
    .Q_N(_0536_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[7] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net63),
    .D(net196),
    .Q_N(_0014_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[0] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net61),
    .D(_0043_),
    .Q_N(_0535_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net59),
    .D(_0044_),
    .Q_N(_0008_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[2] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net57),
    .D(_0045_),
    .Q_N(_0534_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[0] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net55),
    .D(_0046_),
    .Q_N(_0533_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[1] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net53),
    .D(_0047_),
    .Q_N(_0532_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[2] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net51),
    .D(_0048_),
    .Q_N(_0531_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[3] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net49),
    .D(_0049_),
    .Q_N(_0530_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[4] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net47),
    .D(net268),
    .Q_N(_0529_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[5] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net45),
    .D(_0051_),
    .Q_N(_0528_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[6] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net41),
    .D(_0052_),
    .Q_N(_0527_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[7] ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net39),
    .D(_0053_),
    .Q_N(_0526_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[8] ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net37),
    .D(_0054_),
    .Q_N(_0525_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[9] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net35),
    .D(_0055_),
    .Q_N(_0524_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[10] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net33),
    .D(net297),
    .Q_N(_0523_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[11] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net31),
    .D(_0057_),
    .Q_N(_0522_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[12] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net29),
    .D(net275),
    .Q_N(_0521_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[13] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net27),
    .D(_0059_),
    .Q_N(_0520_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[14] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net25),
    .D(_0060_),
    .Q_N(_0519_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[15] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net23),
    .D(_0061_),
    .Q_N(_0518_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[16] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net164),
    .D(_0062_),
    .Q_N(_0517_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[17] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net162),
    .D(_0063_),
    .Q_N(_0516_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[18] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net160),
    .D(_0064_),
    .Q_N(_0515_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[19] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net158),
    .D(_0065_),
    .Q_N(_0514_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[20] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net156),
    .D(net260),
    .Q_N(_0513_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[21] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net154),
    .D(_0067_),
    .Q_N(_0512_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[22] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net152),
    .D(_0068_),
    .Q_N(_0511_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[23] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net150),
    .D(net218),
    .Q_N(_0510_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[24] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net148),
    .D(_0070_),
    .Q_N(_0509_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[25] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net146),
    .D(net216),
    .Q_N(_0508_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[26] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0072_),
    .Q_N(_0507_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[27] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net142),
    .D(_0073_),
    .Q_N(_0506_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[28] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net140),
    .D(_0074_),
    .Q_N(_0505_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[29] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net138),
    .D(_0075_),
    .Q_N(_0504_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[30] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net136),
    .D(_0076_),
    .Q_N(_0503_),
    .Q(\TRNG_inst.U3_Main_controller.tmp_reg[31] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net134),
    .D(net203),
    .Q_N(_0502_),
    .Q(\TRNG_inst.TX_Active ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net133),
    .D(_0078_),
    .Q_N(_0501_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_RX_DV ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net132),
    .D(_0079_),
    .Q_N(_0013_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[0] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(net378),
    .Q_N(_0500_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[1] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net128),
    .D(net251),
    .Q_N(_0499_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[2] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net126),
    .D(net312),
    .Q_N(_0498_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[3] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net124),
    .D(net272),
    .Q_N(_0497_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[4] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net122),
    .D(net309),
    .Q_N(_0496_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[5] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net91),
    .D(_0085_),
    .Q_N(_0495_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[6] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net62),
    .D(net223),
    .Q_N(_0494_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[7] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net58),
    .D(net317),
    .Q_N(_0493_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[8] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net54),
    .D(_0088_),
    .Q_N(_0492_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[9] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net50),
    .D(net258),
    .Q_N(_0491_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_delay[10] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net46),
    .D(_0090_),
    .Q_N(_0001_),
    .Q(\TRNG_inst.U3_Main_controller.state[2] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net40),
    .D(_0091_),
    .Q_N(_0490_),
    .Q(\TRNG_inst.U3_Main_controller.state[1] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net36),
    .D(net392),
    .Q_N(_0489_),
    .Q(\TRNG_inst.U3_Main_controller.state[0] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net32),
    .D(net329),
    .Q_N(_0488_),
    .Q(\TRNG_inst.TX_Serial ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net28),
    .D(_0094_),
    .Q_N(_0000_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[2] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net26),
    .D(net390),
    .Q_N(_0487_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[1] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net24),
    .D(net382),
    .Q_N(_0486_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[0] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net165),
    .D(net344),
    .Q_N(_0485_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[9] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net161),
    .D(net307),
    .Q_N(_0004_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[8] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net157),
    .D(net323),
    .Q_N(_0005_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net153),
    .D(net342),
    .Q_N(_0007_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net149),
    .D(net331),
    .Q_N(_0484_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(net326),
    .Q_N(_0483_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[4] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net141),
    .D(net354),
    .Q_N(_0006_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[3] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net137),
    .D(net356),
    .Q_N(_0482_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net131),
    .D(net320),
    .Q_N(_0481_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[1] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net127),
    .D(_0106_),
    .Q_N(_0480_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net123),
    .D(net351),
    .Q_N(_0003_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[2] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net121),
    .D(net337),
    .Q_N(_0479_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[1] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net90),
    .D(net373),
    .Q_N(_0478_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net60),
    .D(net371),
    .Q_N(_0477_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net52),
    .D(_0111_),
    .Q_N(_0476_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[8] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net44),
    .D(net303),
    .Q_N(_0475_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[7] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net34),
    .D(_0113_),
    .Q_N(_0474_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[6] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net163),
    .D(_0114_),
    .Q_N(_0473_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net155),
    .D(_0115_),
    .Q_N(_0472_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[4] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net147),
    .D(_0116_),
    .Q_N(_0471_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[3] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net139),
    .D(_0117_),
    .Q_N(_0470_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net129),
    .D(_0118_),
    .Q_N(_0469_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net56),
    .D(_0119_),
    .Q_N(_0468_),
    .Q(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[0] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net38),
    .D(net205),
    .Q_N(_0467_),
    .Q(\TRNG_inst.TX_DV ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net159),
    .D(net193),
    .Q_N(_0012_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[0] ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net143),
    .D(net340),
    .Q_N(_0466_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net125),
    .D(net348),
    .Q_N(_0002_),
    .Q(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[2] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net30),
    .D(net188),
    .Q_N(_0011_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_bytes[0] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net135),
    .D(net365),
    .Q_N(_0465_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_bytes[1] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net151),
    .D(_0126_),
    .Q_N(_0010_),
    .Q(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ));
 sg13g2_tiehi _1211__24 (.L_HI(net24));
 sg13g2_tiehi _1175__25 (.L_HI(net25));
 sg13g2_tiehi _1210__26 (.L_HI(net26));
 sg13g2_tiehi _1174__27 (.L_HI(net27));
 sg13g2_tiehi _1209__28 (.L_HI(net28));
 sg13g2_tiehi _1173__29 (.L_HI(net29));
 sg13g2_tiehi _1239__30 (.L_HI(net30));
 sg13g2_tiehi _1172__31 (.L_HI(net31));
 sg13g2_tiehi _1208__32 (.L_HI(net32));
 sg13g2_tiehi _1171__33 (.L_HI(net33));
 sg13g2_tiehi _1228__34 (.L_HI(net34));
 sg13g2_tiehi _1170__35 (.L_HI(net35));
 sg13g2_tiehi _1207__36 (.L_HI(net36));
 sg13g2_tiehi _1169__37 (.L_HI(net37));
 sg13g2_tiehi _1235__38 (.L_HI(net38));
 sg13g2_tiehi _1168__39 (.L_HI(net39));
 sg13g2_tiehi _1206__40 (.L_HI(net40));
 sg13g2_tiehi _1167__41 (.L_HI(net41));
 sg13g2_tiehi _1128__42 (.L_HI(net42));
 sg13g2_tiehi _1146__43 (.L_HI(net43));
 sg13g2_tiehi _1227__44 (.L_HI(net44));
 sg13g2_tiehi _1166__45 (.L_HI(net45));
 sg13g2_tiehi _1205__46 (.L_HI(net46));
 sg13g2_tiehi _1165__47 (.L_HI(net47));
 sg13g2_tiehi _1147__48 (.L_HI(net48));
 sg13g2_tiehi _1164__49 (.L_HI(net49));
 sg13g2_tiehi _1204__50 (.L_HI(net50));
 sg13g2_tiehi _1163__51 (.L_HI(net51));
 sg13g2_tiehi _1226__52 (.L_HI(net52));
 sg13g2_tiehi _1162__53 (.L_HI(net53));
 sg13g2_tiehi _1203__54 (.L_HI(net54));
 sg13g2_tiehi _1161__55 (.L_HI(net55));
 sg13g2_tiehi _1234__56 (.L_HI(net56));
 sg13g2_tiehi _1160__57 (.L_HI(net57));
 sg13g2_tiehi _1202__58 (.L_HI(net58));
 sg13g2_tiehi _1159__59 (.L_HI(net59));
 sg13g2_tiehi _1225__60 (.L_HI(net60));
 sg13g2_tiehi _1158__61 (.L_HI(net61));
 sg13g2_tiehi _1201__62 (.L_HI(net62));
 sg13g2_tiehi _1157__63 (.L_HI(net63));
 sg13g2_tiehi _1156__64 (.L_HI(net64));
 sg13g2_tiehi _1155__65 (.L_HI(net65));
 sg13g2_tiehi _1154__66 (.L_HI(net66));
 sg13g2_tiehi _1153__67 (.L_HI(net67));
 sg13g2_tiehi _1152__68 (.L_HI(net68));
 sg13g2_tiehi _1151__69 (.L_HI(net69));
 sg13g2_tiehi _1150__70 (.L_HI(net70));
 sg13g2_tiehi _1149__71 (.L_HI(net71));
 sg13g2_tiehi _1148__72 (.L_HI(net72));
 sg13g2_tiehi _1145__73 (.L_HI(net73));
 sg13g2_tiehi _1144__74 (.L_HI(net74));
 sg13g2_tiehi _1143__75 (.L_HI(net75));
 sg13g2_tiehi _1142__76 (.L_HI(net76));
 sg13g2_tiehi _1141__77 (.L_HI(net77));
 sg13g2_tiehi _1140__78 (.L_HI(net78));
 sg13g2_tiehi _1139__79 (.L_HI(net79));
 sg13g2_tiehi _1138__80 (.L_HI(net80));
 sg13g2_tiehi _1137__81 (.L_HI(net81));
 sg13g2_tiehi _1136__82 (.L_HI(net82));
 sg13g2_tiehi _1135__83 (.L_HI(net83));
 sg13g2_tiehi _1134__84 (.L_HI(net84));
 sg13g2_tiehi _1133__85 (.L_HI(net85));
 sg13g2_tiehi _1132__86 (.L_HI(net86));
 sg13g2_tiehi _1131__87 (.L_HI(net87));
 sg13g2_tiehi _1130__88 (.L_HI(net88));
 sg13g2_tiehi _1129__89 (.L_HI(net89));
 sg13g2_tiehi _1224__90 (.L_HI(net90));
 sg13g2_tiehi _1200__91 (.L_HI(net91));
 sg13g2_tiehi _1223__92 (.L_HI(net121));
 sg13g2_tiehi _1199__93 (.L_HI(net122));
 sg13g2_tiehi _1222__94 (.L_HI(net123));
 sg13g2_tiehi _1198__95 (.L_HI(net124));
 sg13g2_tiehi _1238__96 (.L_HI(net125));
 sg13g2_tiehi _1197__97 (.L_HI(net126));
 sg13g2_tiehi _1221__98 (.L_HI(net127));
 sg13g2_tiehi _1196__99 (.L_HI(net128));
 sg13g2_tiehi _1233__100 (.L_HI(net129));
 sg13g2_tiehi _1195__101 (.L_HI(net130));
 sg13g2_tiehi _1220__102 (.L_HI(net131));
 sg13g2_tiehi _1194__103 (.L_HI(net132));
 sg13g2_tiehi _1193__104 (.L_HI(net133));
 sg13g2_tiehi _1192__105 (.L_HI(net134));
 sg13g2_tiehi _1240__106 (.L_HI(net135));
 sg13g2_tiehi _1191__107 (.L_HI(net136));
 sg13g2_tiehi _1219__108 (.L_HI(net137));
 sg13g2_tiehi _1190__109 (.L_HI(net138));
 sg13g2_tiehi _1232__110 (.L_HI(net139));
 sg13g2_tiehi _1189__111 (.L_HI(net140));
 sg13g2_tiehi _1218__112 (.L_HI(net141));
 sg13g2_tiehi _1188__113 (.L_HI(net142));
 sg13g2_tiehi _1237__114 (.L_HI(net143));
 sg13g2_tiehi _1187__115 (.L_HI(net144));
 sg13g2_tiehi _1217__116 (.L_HI(net145));
 sg13g2_tiehi _1186__117 (.L_HI(net146));
 sg13g2_tiehi _1231__118 (.L_HI(net147));
 sg13g2_tiehi _1185__119 (.L_HI(net148));
 sg13g2_tiehi _1216__120 (.L_HI(net149));
 sg13g2_tiehi _1184__121 (.L_HI(net150));
 sg13g2_tiehi _1241__122 (.L_HI(net151));
 sg13g2_tiehi _1183__123 (.L_HI(net152));
 sg13g2_tiehi _1215__124 (.L_HI(net153));
 sg13g2_tiehi _1182__125 (.L_HI(net154));
 sg13g2_tiehi _1230__126 (.L_HI(net155));
 sg13g2_tiehi _1181__127 (.L_HI(net156));
 sg13g2_tiehi _1214__128 (.L_HI(net157));
 sg13g2_tiehi _1180__129 (.L_HI(net158));
 sg13g2_tiehi _1236__130 (.L_HI(net159));
 sg13g2_tiehi _1179__131 (.L_HI(net160));
 sg13g2_tiehi _1213__132 (.L_HI(net161));
 sg13g2_tiehi _1178__133 (.L_HI(net162));
 sg13g2_tiehi _1229__134 (.L_HI(net163));
 sg13g2_tiehi _1177__135 (.L_HI(net164));
 sg13g2_tiehi _1212__136 (.L_HI(net165));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_daobaanh_rng_4 (.L_LO(net4));
 sg13g2_tielo tt_um_daobaanh_rng_5 (.L_LO(net5));
 sg13g2_tielo tt_um_daobaanh_rng_6 (.L_LO(net6));
 sg13g2_tielo tt_um_daobaanh_rng_7 (.L_LO(net7));
 sg13g2_tielo tt_um_daobaanh_rng_8 (.L_LO(net8));
 sg13g2_tielo tt_um_daobaanh_rng_9 (.L_LO(net9));
 sg13g2_tielo tt_um_daobaanh_rng_10 (.L_LO(net10));
 sg13g2_tielo tt_um_daobaanh_rng_11 (.L_LO(net11));
 sg13g2_tielo tt_um_daobaanh_rng_12 (.L_LO(net12));
 sg13g2_tielo tt_um_daobaanh_rng_13 (.L_LO(net13));
 sg13g2_tielo tt_um_daobaanh_rng_14 (.L_LO(net14));
 sg13g2_tielo tt_um_daobaanh_rng_15 (.L_LO(net15));
 sg13g2_tielo tt_um_daobaanh_rng_16 (.L_LO(net16));
 sg13g2_tielo tt_um_daobaanh_rng_17 (.L_LO(net17));
 sg13g2_tielo tt_um_daobaanh_rng_18 (.L_LO(net18));
 sg13g2_tielo tt_um_daobaanh_rng_19 (.L_LO(net19));
 sg13g2_tielo tt_um_daobaanh_rng_20 (.L_LO(net20));
 sg13g2_tielo tt_um_daobaanh_rng_21 (.L_LO(net21));
 sg13g2_tielo tt_um_daobaanh_rng_22 (.L_LO(net22));
 sg13g2_tiehi _1176__23 (.L_HI(net23));
 sg13g2_buf_2 _1376_ (.A(\TRNG_inst.TX_Serial ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1377_ (.A(\TRNG_inst.U1_TRNG.o_RNG ),
    .X(uo_out[2]));
 sg13g2_buf_2 _1378_ (.A(\TRNG_inst.U3_Main_controller.led ),
    .X(uo_out[3]));
 sg13g2_buf_2 fanout92 (.A(_0377_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net95),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0290_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0215_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net102),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(net104),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0291_),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_0239_));
 sg13g2_buf_2 fanout106 (.A(net108),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0209_),
    .X(net108));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(_0205_));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_0203_));
 sg13g2_buf_2 fanout111 (.A(_0003_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net324),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net387),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(net386));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net386),
    .X(net120));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_tielo tt_um_daobaanh_rng_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Data_R ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold2 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[22] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold3 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold4 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[13] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold5 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[24] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold6 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[18] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold7 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[19] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold8 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[21] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold9 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[11] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold10 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[9] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold11 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[26] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold12 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[27] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold13 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[15] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold14 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[30] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold15 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[16] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold16 (.A(\TRNG_inst.U1_TRNG.o_RNG ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold17 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold18 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[29] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold19 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[7] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold20 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0011_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0459_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0124_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0013_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0328_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0012_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0452_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0121_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold29 (.A(\TRNG_inst.U1_TRNG.o_data[7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0014_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0042_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold32 (.A(\TRNG_inst.U1_TRNG.o_data[9] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold33 (.A(\TRNG_inst.U1_TRNG.o_data[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold34 (.A(\TRNG_inst.U1_TRNG.o_data[29] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold35 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[7] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold36 (.A(\TRNG_inst.U1_TRNG.o_data[15] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold37 (.A(\TRNG_inst.TX_Active ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0077_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold39 (.A(\TRNG_inst.TX_DV ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0120_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold41 (.A(\TRNG_inst.U1_TRNG.o_data[1] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold42 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0015_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold44 (.A(\TRNG_inst.TX_Byte[7] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0033_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold46 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0251_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0034_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold49 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold50 (.A(\TRNG_inst.U1_TRNG.o_data[26] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0071_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold52 (.A(\TRNG_inst.U1_TRNG.o_data[24] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0069_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold54 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[5] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0039_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold56 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[3] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold57 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[7] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0086_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold59 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[9] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold60 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0260_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0036_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold63 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[29] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold64 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[15] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold65 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[23] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0237_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold67 (.A(\TRNG_inst.TX_Byte[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0019_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold69 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[28] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold70 (.A(\TRNG_inst.U1_TRNG.o_data[18] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold71 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[17] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold72 (.A(\TRNG_inst.TX_Byte[4] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0022_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold74 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0267_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0038_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold77 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[16] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold78 (.A(\TRNG_inst.TX_Byte[0] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0018_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold80 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[8] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold81 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[22] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold82 (.A(\TRNG_inst.TX_Byte[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0024_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold84 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[31] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold85 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[2] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0081_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold87 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[30] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold88 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[25] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold89 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[18] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold90 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[7] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0041_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold92 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[10] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0089_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold94 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[21] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0066_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold96 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold97 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[17] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold98 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[10] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold99 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold100 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[1] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0035_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold102 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0050_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold104 (.A(\TRNG_inst.U3_Main_controller.led ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0016_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold106 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[4] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0083_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold108 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[12] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold109 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[13] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0058_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold111 (.A(\TRNG_inst.TX_Byte[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0020_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold113 (.A(\TRNG_inst.U1_TRNG.o_data[21] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold114 (.A(\TRNG_inst.U1_TRNG.RG_part/i_r[20] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold115 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0442_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold117 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[6] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold118 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[4] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold119 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold120 (.A(\TRNG_inst.TX_Byte[3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0021_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold122 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[19] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold123 (.A(\TRNG_inst.TX_Byte[5] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold124 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[2] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold125 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[27] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold126 (.A(\TRNG_inst.U1_TRNG.o_data[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold127 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[6] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0271_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0040_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold130 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold131 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[11] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0056_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold133 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[20] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold134 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_RX_Byte[3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0037_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold136 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[14] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold137 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[7] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0112_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold139 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[5] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold140 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_TX_Data[3] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold141 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[8] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0098_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold143 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[5] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0084_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold145 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[0] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold146 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[3] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0082_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold148 (.A(\TRNG_inst.U3_Main_controller.tmp_reg[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold149 (.A(\TRNG_inst.U1_TRNG.o_data[11] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold150 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold151 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[8] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0087_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold153 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0400_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0105_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold156 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[4] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold157 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[7] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0099_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0000_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0394_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0102_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold162 (.A(\TRNG_inst.TX_Serial ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0359_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0093_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold165 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[5] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0101_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold167 (.A(\TRNG_inst.U1_TRNG.o_data[13] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold168 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[8] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0429_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold170 (.A(\TRNG_inst.U3_Main_controller.state[2] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0009_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0108_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold173 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[1] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0454_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0122_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold176 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0100_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold178 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[9] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0097_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold180 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold181 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[0] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold182 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Bit_Index[2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0123_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold184 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0246_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0107_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0006_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0397_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0103_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold190 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_Clk_Count[2] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0104_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold192 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[2] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0326_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0327_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0001_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0198_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0017_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold198 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[5] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold199 (.A(\TRNG_inst.U3_Main_controller.cnt_bytes[1] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0125_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold201 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold202 (.A(\TRNG_inst.U3_Main_controller.cnt_bytes[2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0464_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold204 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[2] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold205 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[9] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0110_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold207 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_SM_Main[0] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0109_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold209 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[9] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold210 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[6] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold211 (.A(\TRNG_inst.U3_Main_controller.cnt_delay[1] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0330_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0080_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold214 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Clk_Count[6] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold215 (.A(\TRNG_inst.U2_UART_interface.RX_part.r_Bit_Index[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0002_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0096_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold218 (.A(\TRNG_inst.U2_UART_interface.TX_part.r_SM_Main[1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0191_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0192_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold221 (.A(\TRNG_inst.U1_TRNG.i_rst ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold222 (.A(\TRNG_inst.U3_Main_controller.state[1] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0346_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0005_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0095_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold226 (.A(\TRNG_inst.U3_Main_controller.state[0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0092_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0001_),
    .X(net393));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_139 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_4 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_197 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_fill_2 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_decap_4 FILLER_10_160 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_4 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_302 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_324 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_370 ();
 sg13g2_fill_2 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_4 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_decap_4 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_4 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_fill_1 FILLER_11_345 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_fill_2 FILLER_11_391 ();
 sg13g2_fill_1 FILLER_11_393 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_117 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_4 FILLER_13_284 ();
 sg13g2_decap_4 FILLER_13_292 ();
 sg13g2_fill_2 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_355 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_4 FILLER_15_255 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_fill_2 FILLER_15_390 ();
 sg13g2_fill_1 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_86 ();
 sg13g2_decap_8 FILLER_16_93 ();
 sg13g2_decap_8 FILLER_16_100 ();
 sg13g2_decap_4 FILLER_16_107 ();
 sg13g2_fill_1 FILLER_16_111 ();
 sg13g2_fill_2 FILLER_16_162 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_2 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_306 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_49 ();
 sg13g2_decap_4 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_decap_4 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_331 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_4 FILLER_18_25 ();
 sg13g2_fill_1 FILLER_18_29 ();
 sg13g2_fill_2 FILLER_18_33 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_268 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_decap_4 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_243 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_59 ();
 sg13g2_decap_8 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_87 ();
 sg13g2_decap_4 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_145 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_16 ();
 sg13g2_fill_1 FILLER_21_18 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_2 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_fill_1 FILLER_23_50 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_16 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_decap_4 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_11 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_decap_4 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_decap_4 FILLER_28_120 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_4 FILLER_28_138 ();
 sg13g2_fill_2 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_11 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_69 ();
 sg13g2_decap_4 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_37 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_64 ();
 sg13g2_fill_1 FILLER_32_66 ();
 sg13g2_decap_4 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_fill_2 FILLER_32_341 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_22 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_82 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_72 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_decap_8 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_2 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_106 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_257 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_399 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[4] = net19;
 assign uo_out[5] = net20;
 assign uo_out[6] = net21;
 assign uo_out[7] = net22;
endmodule

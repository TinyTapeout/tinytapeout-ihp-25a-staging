module tt_um_i2s_to_pwm_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire \u_top_module.i2s_data_L[10] ;
 wire \u_top_module.i2s_data_L[11] ;
 wire \u_top_module.i2s_data_L[12] ;
 wire \u_top_module.i2s_data_L[13] ;
 wire \u_top_module.i2s_data_L[14] ;
 wire \u_top_module.i2s_data_L[15] ;
 wire \u_top_module.i2s_data_L[8] ;
 wire \u_top_module.i2s_data_L[9] ;
 wire \u_top_module.i2s_data_R[10] ;
 wire \u_top_module.i2s_data_R[11] ;
 wire \u_top_module.i2s_data_R[12] ;
 wire \u_top_module.i2s_data_R[13] ;
 wire \u_top_module.i2s_data_R[14] ;
 wire \u_top_module.i2s_data_R[15] ;
 wire \u_top_module.i2s_data_R[8] ;
 wire \u_top_module.i2s_data_R[9] ;
 wire \u_top_module.left_channel ;
 wire \u_top_module.right_channel ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[0] ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[1] ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[2] ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[3] ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[4] ;
 wire \u_top_module.u_i2s_rx_64x.bit_count[5] ;
 wire \u_top_module.u_i2s_rx_64x.lrclk_prev ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[0] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[10] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[11] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[12] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[13] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[14] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[15] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[1] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[2] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[3] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[4] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[5] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[6] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[7] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[8] ;
 wire \u_top_module.u_i2s_rx_64x.shift_reg[9] ;
 wire \u_top_module.u_pwm_generator_L.counter[0] ;
 wire \u_top_module.u_pwm_generator_L.counter[1] ;
 wire \u_top_module.u_pwm_generator_L.counter[2] ;
 wire \u_top_module.u_pwm_generator_L.counter[3] ;
 wire \u_top_module.u_pwm_generator_L.counter[4] ;
 wire \u_top_module.u_pwm_generator_L.counter[5] ;
 wire \u_top_module.u_pwm_generator_L.counter[6] ;
 wire \u_top_module.u_pwm_generator_L.counter[7] ;
 wire \u_top_module.u_pwm_generator_R.counter[0] ;
 wire \u_top_module.u_pwm_generator_R.counter[1] ;
 wire \u_top_module.u_pwm_generator_R.counter[2] ;
 wire \u_top_module.u_pwm_generator_R.counter[3] ;
 wire \u_top_module.u_pwm_generator_R.counter[4] ;
 wire \u_top_module.u_pwm_generator_R.counter[5] ;
 wire \u_top_module.u_pwm_generator_R.counter[6] ;
 wire \u_top_module.u_pwm_generator_R.counter[7] ;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;

 sg13g2_inv_1 _198_ (.Y(_056_),
    .A(\u_top_module.u_pwm_generator_L.counter[5] ));
 sg13g2_inv_1 _199_ (.Y(_057_),
    .A(\u_top_module.i2s_data_L[11] ));
 sg13g2_inv_1 _200_ (.Y(_058_),
    .A(\u_top_module.u_pwm_generator_L.counter[3] ));
 sg13g2_inv_1 _201_ (.Y(_059_),
    .A(\u_top_module.u_pwm_generator_L.counter[2] ));
 sg13g2_inv_1 _202_ (.Y(_060_),
    .A(\u_top_module.u_pwm_generator_L.counter[1] ));
 sg13g2_inv_1 _203_ (.Y(_006_),
    .A(\u_top_module.u_pwm_generator_L.counter[0] ));
 sg13g2_inv_1 _204_ (.Y(_015_),
    .A(\u_top_module.u_pwm_generator_R.counter[0] ));
 sg13g2_inv_1 _205_ (.Y(_061_),
    .A(\u_top_module.u_pwm_generator_R.counter[3] ));
 sg13g2_inv_1 _206_ (.Y(_062_),
    .A(\u_top_module.u_pwm_generator_R.counter[6] ));
 sg13g2_inv_1 _207_ (.Y(_063_),
    .A(\u_top_module.u_pwm_generator_R.counter[7] ));
 sg13g2_inv_1 _208_ (.Y(_064_),
    .A(\u_top_module.u_pwm_generator_L.counter[7] ));
 sg13g2_inv_1 _209_ (.Y(_065_),
    .A(\u_top_module.i2s_data_R[13] ));
 sg13g2_nand2_1 _210_ (.Y(_066_),
    .A(_064_),
    .B(\u_top_module.i2s_data_L[15] ));
 sg13g2_nand2b_1 _211_ (.Y(_067_),
    .B(\u_top_module.u_pwm_generator_L.counter[4] ),
    .A_N(\u_top_module.i2s_data_L[12] ));
 sg13g2_o21ai_1 _212_ (.B1(_067_),
    .Y(_068_),
    .A1(\u_top_module.i2s_data_L[13] ),
    .A2(_056_));
 sg13g2_nand2_1 _213_ (.Y(_069_),
    .A(\u_top_module.i2s_data_L[13] ),
    .B(_056_));
 sg13g2_nand2b_1 _214_ (.Y(_070_),
    .B(\u_top_module.i2s_data_L[14] ),
    .A_N(\u_top_module.u_pwm_generator_L.counter[6] ));
 sg13g2_nand3_1 _215_ (.B(_069_),
    .C(_070_),
    .A(_068_),
    .Y(_071_));
 sg13g2_nand2b_1 _216_ (.Y(_072_),
    .B(\u_top_module.u_pwm_generator_L.counter[6] ),
    .A_N(\u_top_module.i2s_data_L[14] ));
 sg13g2_o21ai_1 _217_ (.B1(_072_),
    .Y(_073_),
    .A1(_064_),
    .A2(\u_top_module.i2s_data_L[15] ));
 sg13g2_nand2b_1 _218_ (.Y(_074_),
    .B(_071_),
    .A_N(_073_));
 sg13g2_nand2b_1 _219_ (.Y(_075_),
    .B(\u_top_module.u_pwm_generator_L.counter[1] ),
    .A_N(\u_top_module.i2s_data_L[9] ));
 sg13g2_nand3_1 _220_ (.B(_006_),
    .C(_075_),
    .A(\u_top_module.i2s_data_L[8] ),
    .Y(_076_));
 sg13g2_a22oi_1 _221_ (.Y(_077_),
    .B1(\u_top_module.i2s_data_L[9] ),
    .B2(_060_),
    .A2(_059_),
    .A1(\u_top_module.i2s_data_L[10] ));
 sg13g2_nor2_1 _222_ (.A(\u_top_module.i2s_data_L[10] ),
    .B(_059_),
    .Y(_078_));
 sg13g2_a221oi_1 _223_ (.B2(_077_),
    .C1(_078_),
    .B1(_076_),
    .A1(_057_),
    .Y(_079_),
    .A2(\u_top_module.u_pwm_generator_L.counter[3] ));
 sg13g2_nand2b_1 _224_ (.Y(_080_),
    .B(\u_top_module.i2s_data_L[12] ),
    .A_N(\u_top_module.u_pwm_generator_L.counter[4] ));
 sg13g2_nand4_1 _225_ (.B(_070_),
    .C(_072_),
    .A(_069_),
    .Y(_081_),
    .D(_080_));
 sg13g2_o21ai_1 _226_ (.B1(_066_),
    .Y(_082_),
    .A1(_057_),
    .A2(\u_top_module.u_pwm_generator_L.counter[3] ));
 sg13g2_nor4_1 _227_ (.A(_068_),
    .B(_079_),
    .C(_081_),
    .D(_082_),
    .Y(_083_));
 sg13g2_a21oi_1 _228_ (.A1(_066_),
    .A2(_074_),
    .Y(_014_),
    .B1(_083_));
 sg13g2_xor2_1 _229_ (.B(\u_top_module.u_pwm_generator_R.counter[0] ),
    .A(\u_top_module.u_pwm_generator_R.counter[1] ),
    .X(_016_));
 sg13g2_nand3_1 _230_ (.B(\u_top_module.u_pwm_generator_R.counter[0] ),
    .C(\u_top_module.u_pwm_generator_R.counter[2] ),
    .A(\u_top_module.u_pwm_generator_R.counter[1] ),
    .Y(_084_));
 sg13g2_a21o_1 _231_ (.A2(\u_top_module.u_pwm_generator_R.counter[0] ),
    .A1(\u_top_module.u_pwm_generator_R.counter[1] ),
    .B1(\u_top_module.u_pwm_generator_R.counter[2] ),
    .X(_085_));
 sg13g2_and2_1 _232_ (.A(_084_),
    .B(_085_),
    .X(_017_));
 sg13g2_nor2_1 _233_ (.A(_061_),
    .B(_084_),
    .Y(_086_));
 sg13g2_xnor2_1 _234_ (.Y(_018_),
    .A(\u_top_module.u_pwm_generator_R.counter[3] ),
    .B(_084_));
 sg13g2_xor2_1 _235_ (.B(_086_),
    .A(\u_top_module.u_pwm_generator_R.counter[4] ),
    .X(_019_));
 sg13g2_nand3_1 _236_ (.B(\u_top_module.u_pwm_generator_R.counter[4] ),
    .C(_086_),
    .A(\u_top_module.u_pwm_generator_R.counter[5] ),
    .Y(_087_));
 sg13g2_a21o_1 _237_ (.A2(_086_),
    .A1(\u_top_module.u_pwm_generator_R.counter[4] ),
    .B1(\u_top_module.u_pwm_generator_R.counter[5] ),
    .X(_088_));
 sg13g2_and2_1 _238_ (.A(_087_),
    .B(_088_),
    .X(_020_));
 sg13g2_or2_1 _239_ (.X(_089_),
    .B(_087_),
    .A(_063_));
 sg13g2_xnor2_1 _240_ (.Y(_090_),
    .A(\u_top_module.u_pwm_generator_R.counter[6] ),
    .B(_087_));
 sg13g2_and2_1 _241_ (.A(_089_),
    .B(_090_),
    .X(_021_));
 sg13g2_o21ai_1 _242_ (.B1(_063_),
    .Y(_091_),
    .A1(_062_),
    .A2(_087_));
 sg13g2_and2_1 _243_ (.A(_089_),
    .B(_091_),
    .X(_022_));
 sg13g2_xor2_1 _244_ (.B(\u_top_module.u_pwm_generator_L.counter[0] ),
    .A(\u_top_module.u_pwm_generator_L.counter[1] ),
    .X(_007_));
 sg13g2_nand3_1 _245_ (.B(\u_top_module.u_pwm_generator_L.counter[1] ),
    .C(\u_top_module.u_pwm_generator_L.counter[0] ),
    .A(\u_top_module.u_pwm_generator_L.counter[2] ),
    .Y(_092_));
 sg13g2_o21ai_1 _246_ (.B1(_059_),
    .Y(_093_),
    .A1(_060_),
    .A2(_006_));
 sg13g2_and2_1 _247_ (.A(_092_),
    .B(_093_),
    .X(_008_));
 sg13g2_nor2_1 _248_ (.A(_058_),
    .B(_092_),
    .Y(_094_));
 sg13g2_xnor2_1 _249_ (.Y(_009_),
    .A(\u_top_module.u_pwm_generator_L.counter[3] ),
    .B(_092_));
 sg13g2_xor2_1 _250_ (.B(_094_),
    .A(\u_top_module.u_pwm_generator_L.counter[4] ),
    .X(_010_));
 sg13g2_and3_1 _251_ (.X(_095_),
    .A(\u_top_module.u_pwm_generator_L.counter[5] ),
    .B(\u_top_module.u_pwm_generator_L.counter[4] ),
    .C(_094_));
 sg13g2_a21oi_1 _252_ (.A1(\u_top_module.u_pwm_generator_L.counter[4] ),
    .A2(_094_),
    .Y(_096_),
    .B1(\u_top_module.u_pwm_generator_L.counter[5] ));
 sg13g2_nor2_1 _253_ (.A(_095_),
    .B(_096_),
    .Y(_011_));
 sg13g2_a21oi_1 _254_ (.A1(_064_),
    .A2(_095_),
    .Y(_097_),
    .B1(\u_top_module.u_pwm_generator_L.counter[6] ));
 sg13g2_a21oi_1 _255_ (.A1(\u_top_module.u_pwm_generator_L.counter[6] ),
    .A2(_095_),
    .Y(_012_),
    .B1(_097_));
 sg13g2_a21oi_1 _256_ (.A1(\u_top_module.u_pwm_generator_L.counter[6] ),
    .A2(_095_),
    .Y(_098_),
    .B1(\u_top_module.u_pwm_generator_L.counter[7] ));
 sg13g2_a21oi_1 _257_ (.A1(\u_top_module.u_pwm_generator_L.counter[7] ),
    .A2(_095_),
    .Y(_013_),
    .B1(_098_));
 sg13g2_nor2b_2 _258_ (.A(net3),
    .B_N(\u_top_module.u_i2s_rx_64x.lrclk_prev ),
    .Y(_099_));
 sg13g2_nor2b_2 _259_ (.A(\u_top_module.u_i2s_rx_64x.lrclk_prev ),
    .B_N(net3),
    .Y(_100_));
 sg13g2_or2_2 _260_ (.X(_101_),
    .B(net8),
    .A(net9));
 sg13g2_nor2_1 _261_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[0] ),
    .B(_101_),
    .Y(_000_));
 sg13g2_nor2_1 _262_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[0] ),
    .B(\u_top_module.u_i2s_rx_64x.bit_count[1] ),
    .Y(_102_));
 sg13g2_and2_1 _263_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[0] ),
    .B(\u_top_module.u_i2s_rx_64x.bit_count[1] ),
    .X(_103_));
 sg13g2_nor3_1 _264_ (.A(_101_),
    .B(_102_),
    .C(_103_),
    .Y(_001_));
 sg13g2_nor2_1 _265_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[2] ),
    .B(_103_),
    .Y(_104_));
 sg13g2_and2_1 _266_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[2] ),
    .B(_103_),
    .X(_105_));
 sg13g2_nor3_1 _267_ (.A(_101_),
    .B(_104_),
    .C(_105_),
    .Y(_002_));
 sg13g2_nor2_1 _268_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[3] ),
    .B(_105_),
    .Y(_106_));
 sg13g2_and3_1 _269_ (.X(_107_),
    .A(\u_top_module.u_i2s_rx_64x.bit_count[2] ),
    .B(\u_top_module.u_i2s_rx_64x.bit_count[3] ),
    .C(_103_));
 sg13g2_nor3_1 _270_ (.A(_101_),
    .B(_106_),
    .C(_107_),
    .Y(_003_));
 sg13g2_nor2_1 _271_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[4] ),
    .B(_107_),
    .Y(_108_));
 sg13g2_and2_1 _272_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[4] ),
    .B(_107_),
    .X(_109_));
 sg13g2_nor3_1 _273_ (.A(_101_),
    .B(_108_),
    .C(_109_),
    .Y(_004_));
 sg13g2_xnor2_1 _274_ (.Y(_110_),
    .A(\u_top_module.u_i2s_rx_64x.bit_count[5] ),
    .B(_109_));
 sg13g2_nor2_1 _275_ (.A(_101_),
    .B(_110_),
    .Y(_005_));
 sg13g2_nand2b_1 _276_ (.Y(_111_),
    .B(\u_top_module.i2s_data_R[15] ),
    .A_N(\u_top_module.u_pwm_generator_R.counter[7] ));
 sg13g2_nand2b_1 _277_ (.Y(_112_),
    .B(\u_top_module.i2s_data_R[14] ),
    .A_N(\u_top_module.u_pwm_generator_R.counter[6] ));
 sg13g2_nand2_1 _278_ (.Y(_113_),
    .A(_111_),
    .B(_112_));
 sg13g2_nand2b_1 _279_ (.Y(_114_),
    .B(\u_top_module.u_pwm_generator_R.counter[7] ),
    .A_N(\u_top_module.i2s_data_R[15] ));
 sg13g2_nand2b_1 _280_ (.Y(_115_),
    .B(\u_top_module.u_pwm_generator_R.counter[6] ),
    .A_N(\u_top_module.i2s_data_R[14] ));
 sg13g2_nor2b_1 _281_ (.A(\u_top_module.i2s_data_R[13] ),
    .B_N(\u_top_module.u_pwm_generator_R.counter[5] ),
    .Y(_116_));
 sg13g2_nand4_1 _282_ (.B(_112_),
    .C(_114_),
    .A(_111_),
    .Y(_117_),
    .D(_115_));
 sg13g2_nor2_1 _283_ (.A(_116_),
    .B(_117_),
    .Y(_118_));
 sg13g2_nand2b_1 _284_ (.Y(_119_),
    .B(\u_top_module.i2s_data_R[12] ),
    .A_N(\u_top_module.u_pwm_generator_R.counter[4] ));
 sg13g2_o21ai_1 _285_ (.B1(_119_),
    .Y(_120_),
    .A1(\u_top_module.u_pwm_generator_R.counter[5] ),
    .A2(_065_));
 sg13g2_nor2b_1 _286_ (.A(\u_top_module.i2s_data_R[12] ),
    .B_N(\u_top_module.u_pwm_generator_R.counter[4] ),
    .Y(_121_));
 sg13g2_nor4_2 _287_ (.A(_116_),
    .B(_117_),
    .C(_120_),
    .Y(_122_),
    .D(_121_));
 sg13g2_nor2b_1 _288_ (.A(\u_top_module.u_pwm_generator_R.counter[2] ),
    .B_N(\u_top_module.i2s_data_R[10] ),
    .Y(_123_));
 sg13g2_nor2b_1 _289_ (.A(\u_top_module.u_pwm_generator_R.counter[3] ),
    .B_N(\u_top_module.i2s_data_R[11] ),
    .Y(_124_));
 sg13g2_nor2_1 _290_ (.A(_123_),
    .B(_124_),
    .Y(_125_));
 sg13g2_nor2b_1 _291_ (.A(\u_top_module.i2s_data_R[10] ),
    .B_N(\u_top_module.u_pwm_generator_R.counter[2] ),
    .Y(_126_));
 sg13g2_nor2b_1 _292_ (.A(\u_top_module.i2s_data_R[11] ),
    .B_N(\u_top_module.u_pwm_generator_R.counter[3] ),
    .Y(_127_));
 sg13g2_or4_1 _293_ (.A(_123_),
    .B(_124_),
    .C(_126_),
    .D(_127_),
    .X(_128_));
 sg13g2_nand2b_1 _294_ (.Y(_129_),
    .B(\u_top_module.i2s_data_R[9] ),
    .A_N(\u_top_module.u_pwm_generator_R.counter[1] ));
 sg13g2_xnor2_1 _295_ (.Y(_130_),
    .A(\u_top_module.u_pwm_generator_R.counter[1] ),
    .B(\u_top_module.i2s_data_R[9] ));
 sg13g2_o21ai_1 _296_ (.B1(_130_),
    .Y(_131_),
    .A1(_015_),
    .A2(\u_top_module.i2s_data_R[8] ));
 sg13g2_a21oi_1 _297_ (.A1(_129_),
    .A2(_131_),
    .Y(_132_),
    .B1(_128_));
 sg13g2_nor2_1 _298_ (.A(_125_),
    .B(_127_),
    .Y(_133_));
 sg13g2_o21ai_1 _299_ (.B1(_122_),
    .Y(_134_),
    .A1(_132_),
    .A2(_133_));
 sg13g2_a22oi_1 _300_ (.Y(_135_),
    .B1(_118_),
    .B2(_120_),
    .A2(_114_),
    .A1(_113_));
 sg13g2_nor2b_1 _301_ (.A(\u_top_module.u_pwm_generator_R.counter[0] ),
    .B_N(\u_top_module.i2s_data_R[8] ),
    .Y(_136_));
 sg13g2_nor3_1 _302_ (.A(_128_),
    .B(_131_),
    .C(_136_),
    .Y(_137_));
 sg13g2_a22oi_1 _303_ (.Y(_023_),
    .B1(_137_),
    .B2(_122_),
    .A2(_135_),
    .A1(_134_));
 sg13g2_or3_1 _304_ (.A(\u_top_module.u_i2s_rx_64x.bit_count[5] ),
    .B(\u_top_module.u_i2s_rx_64x.bit_count[4] ),
    .C(_101_),
    .X(_138_));
 sg13g2_mux2_1 _305_ (.A0(net4),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[0] ),
    .S(net5),
    .X(_024_));
 sg13g2_mux2_1 _306_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[0] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[1] ),
    .S(net5),
    .X(_025_));
 sg13g2_mux2_1 _307_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[1] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[2] ),
    .S(net5),
    .X(_026_));
 sg13g2_mux2_1 _308_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[2] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[3] ),
    .S(net5),
    .X(_027_));
 sg13g2_mux2_1 _309_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[3] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[4] ),
    .S(net6),
    .X(_028_));
 sg13g2_mux2_1 _310_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[4] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[5] ),
    .S(net5),
    .X(_029_));
 sg13g2_mux2_1 _311_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[5] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[6] ),
    .S(net5),
    .X(_030_));
 sg13g2_mux2_1 _312_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[6] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[7] ),
    .S(net5),
    .X(_031_));
 sg13g2_mux2_1 _313_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[7] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[8] ),
    .S(net5),
    .X(_032_));
 sg13g2_mux2_1 _314_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[8] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[9] ),
    .S(net6),
    .X(_033_));
 sg13g2_mux2_1 _315_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[9] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[10] ),
    .S(net6),
    .X(_034_));
 sg13g2_mux2_1 _316_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[10] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[11] ),
    .S(net7),
    .X(_035_));
 sg13g2_mux2_1 _317_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[11] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[12] ),
    .S(net7),
    .X(_036_));
 sg13g2_mux2_1 _318_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[12] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[13] ),
    .S(net7),
    .X(_037_));
 sg13g2_mux2_1 _319_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[13] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[14] ),
    .S(net7),
    .X(_038_));
 sg13g2_mux2_1 _320_ (.A0(\u_top_module.u_i2s_rx_64x.shift_reg[14] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[15] ),
    .S(net7),
    .X(_039_));
 sg13g2_mux2_1 _321_ (.A0(\u_top_module.i2s_data_L[8] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[8] ),
    .S(net9),
    .X(_040_));
 sg13g2_mux2_1 _322_ (.A0(\u_top_module.i2s_data_L[9] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[9] ),
    .S(_099_),
    .X(_041_));
 sg13g2_mux2_1 _323_ (.A0(\u_top_module.i2s_data_L[10] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[10] ),
    .S(_099_),
    .X(_042_));
 sg13g2_nand2_1 _324_ (.Y(_139_),
    .A(\u_top_module.u_i2s_rx_64x.shift_reg[11] ),
    .B(net9));
 sg13g2_o21ai_1 _325_ (.B1(_139_),
    .Y(_043_),
    .A1(_057_),
    .A2(net9));
 sg13g2_mux2_1 _326_ (.A0(\u_top_module.i2s_data_L[12] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[12] ),
    .S(net9),
    .X(_044_));
 sg13g2_mux2_1 _327_ (.A0(\u_top_module.i2s_data_L[13] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[13] ),
    .S(net9),
    .X(_045_));
 sg13g2_mux2_1 _328_ (.A0(\u_top_module.i2s_data_L[14] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[14] ),
    .S(net9),
    .X(_046_));
 sg13g2_mux2_1 _329_ (.A0(\u_top_module.i2s_data_L[15] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[15] ),
    .S(net9),
    .X(_047_));
 sg13g2_mux2_1 _330_ (.A0(\u_top_module.i2s_data_R[8] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[8] ),
    .S(_100_),
    .X(_048_));
 sg13g2_mux2_1 _331_ (.A0(\u_top_module.i2s_data_R[9] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[9] ),
    .S(_100_),
    .X(_049_));
 sg13g2_mux2_1 _332_ (.A0(\u_top_module.i2s_data_R[10] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[10] ),
    .S(net8),
    .X(_050_));
 sg13g2_mux2_1 _333_ (.A0(\u_top_module.i2s_data_R[11] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[11] ),
    .S(net8),
    .X(_051_));
 sg13g2_mux2_1 _334_ (.A0(\u_top_module.i2s_data_R[12] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[12] ),
    .S(net8),
    .X(_052_));
 sg13g2_nand2_1 _335_ (.Y(_140_),
    .A(\u_top_module.u_i2s_rx_64x.shift_reg[13] ),
    .B(net8));
 sg13g2_o21ai_1 _336_ (.B1(_140_),
    .Y(_053_),
    .A1(_065_),
    .A2(net8));
 sg13g2_mux2_1 _337_ (.A0(\u_top_module.i2s_data_R[14] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[14] ),
    .S(net8),
    .X(_054_));
 sg13g2_mux2_1 _338_ (.A0(\u_top_module.i2s_data_R[15] ),
    .A1(\u_top_module.u_i2s_rx_64x.shift_reg[15] ),
    .S(net8),
    .X(_055_));
 sg13g2_dfrbp_1 _339_ (.CLK(net17),
    .RESET_B(net27),
    .D(_024_),
    .Q_N(_172_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[0] ));
 sg13g2_dfrbp_1 _340_ (.CLK(net17),
    .RESET_B(net27),
    .D(_025_),
    .Q_N(_171_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[1] ));
 sg13g2_dfrbp_1 _341_ (.CLK(net17),
    .RESET_B(net27),
    .D(_026_),
    .Q_N(_170_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[2] ));
 sg13g2_dfrbp_1 _342_ (.CLK(net17),
    .RESET_B(net27),
    .D(_027_),
    .Q_N(_169_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[3] ));
 sg13g2_dfrbp_1 _343_ (.CLK(net17),
    .RESET_B(net27),
    .D(_028_),
    .Q_N(_168_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[4] ));
 sg13g2_dfrbp_1 _344_ (.CLK(net17),
    .RESET_B(net27),
    .D(_029_),
    .Q_N(_167_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[5] ));
 sg13g2_dfrbp_1 _345_ (.CLK(net19),
    .RESET_B(net29),
    .D(_030_),
    .Q_N(_166_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[6] ));
 sg13g2_dfrbp_1 _346_ (.CLK(net19),
    .RESET_B(net29),
    .D(_031_),
    .Q_N(_165_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[7] ));
 sg13g2_dfrbp_1 _347_ (.CLK(net18),
    .RESET_B(net28),
    .D(_032_),
    .Q_N(_164_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[8] ));
 sg13g2_dfrbp_1 _348_ (.CLK(net15),
    .RESET_B(net25),
    .D(_033_),
    .Q_N(_163_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[9] ));
 sg13g2_dfrbp_1 _349_ (.CLK(net15),
    .RESET_B(net25),
    .D(_034_),
    .Q_N(_162_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[10] ));
 sg13g2_dfrbp_1 _350_ (.CLK(net12),
    .RESET_B(net22),
    .D(_035_),
    .Q_N(_161_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[11] ));
 sg13g2_dfrbp_1 _351_ (.CLK(net12),
    .RESET_B(net22),
    .D(_036_),
    .Q_N(_160_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[12] ));
 sg13g2_dfrbp_1 _352_ (.CLK(net11),
    .RESET_B(net21),
    .D(_037_),
    .Q_N(_159_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[13] ));
 sg13g2_dfrbp_1 _353_ (.CLK(net11),
    .RESET_B(net21),
    .D(_038_),
    .Q_N(_158_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[14] ));
 sg13g2_dfrbp_1 _354_ (.CLK(net11),
    .RESET_B(net21),
    .D(_039_),
    .Q_N(_173_),
    .Q(\u_top_module.u_i2s_rx_64x.shift_reg[15] ));
 sg13g2_dfrbp_1 _355_ (.CLK(net15),
    .RESET_B(net25),
    .D(_015_),
    .Q_N(_174_),
    .Q(\u_top_module.u_pwm_generator_R.counter[0] ));
 sg13g2_dfrbp_1 _356_ (.CLK(net15),
    .RESET_B(net25),
    .D(_016_),
    .Q_N(_175_),
    .Q(\u_top_module.u_pwm_generator_R.counter[1] ));
 sg13g2_dfrbp_1 _357_ (.CLK(net12),
    .RESET_B(net22),
    .D(_017_),
    .Q_N(_176_),
    .Q(\u_top_module.u_pwm_generator_R.counter[2] ));
 sg13g2_dfrbp_1 _358_ (.CLK(net12),
    .RESET_B(net22),
    .D(_018_),
    .Q_N(_177_),
    .Q(\u_top_module.u_pwm_generator_R.counter[3] ));
 sg13g2_dfrbp_1 _359_ (.CLK(net10),
    .RESET_B(net20),
    .D(_019_),
    .Q_N(_178_),
    .Q(\u_top_module.u_pwm_generator_R.counter[4] ));
 sg13g2_dfrbp_1 _360_ (.CLK(net10),
    .RESET_B(net20),
    .D(_020_),
    .Q_N(_179_),
    .Q(\u_top_module.u_pwm_generator_R.counter[5] ));
 sg13g2_dfrbp_1 _361_ (.CLK(net10),
    .RESET_B(net20),
    .D(_021_),
    .Q_N(_180_),
    .Q(\u_top_module.u_pwm_generator_R.counter[6] ));
 sg13g2_dfrbp_1 _362_ (.CLK(net10),
    .RESET_B(net20),
    .D(_022_),
    .Q_N(_181_),
    .Q(\u_top_module.u_pwm_generator_R.counter[7] ));
 sg13g2_dfrbp_1 _363_ (.CLK(net11),
    .RESET_B(net21),
    .D(_023_),
    .Q_N(_182_),
    .Q(\u_top_module.right_channel ));
 sg13g2_dfrbp_1 _364_ (.CLK(net15),
    .RESET_B(net25),
    .D(_006_),
    .Q_N(_183_),
    .Q(\u_top_module.u_pwm_generator_L.counter[0] ));
 sg13g2_dfrbp_1 _365_ (.CLK(net15),
    .RESET_B(net25),
    .D(_007_),
    .Q_N(_184_),
    .Q(\u_top_module.u_pwm_generator_L.counter[1] ));
 sg13g2_dfrbp_1 _366_ (.CLK(net16),
    .RESET_B(net26),
    .D(_008_),
    .Q_N(_185_),
    .Q(\u_top_module.u_pwm_generator_L.counter[2] ));
 sg13g2_dfrbp_1 _367_ (.CLK(net16),
    .RESET_B(net26),
    .D(_009_),
    .Q_N(_186_),
    .Q(\u_top_module.u_pwm_generator_L.counter[3] ));
 sg13g2_dfrbp_1 _368_ (.CLK(net12),
    .RESET_B(net22),
    .D(_010_),
    .Q_N(_187_),
    .Q(\u_top_module.u_pwm_generator_L.counter[4] ));
 sg13g2_dfrbp_1 _369_ (.CLK(net12),
    .RESET_B(net22),
    .D(_011_),
    .Q_N(_188_),
    .Q(\u_top_module.u_pwm_generator_L.counter[5] ));
 sg13g2_dfrbp_1 _370_ (.CLK(net13),
    .RESET_B(net23),
    .D(_012_),
    .Q_N(_189_),
    .Q(\u_top_module.u_pwm_generator_L.counter[6] ));
 sg13g2_dfrbp_1 _371_ (.CLK(net13),
    .RESET_B(net23),
    .D(_013_),
    .Q_N(_190_),
    .Q(\u_top_module.u_pwm_generator_L.counter[7] ));
 sg13g2_dfrbp_1 _372_ (.CLK(net11),
    .RESET_B(net21),
    .D(_014_),
    .Q_N(_191_),
    .Q(\u_top_module.left_channel ));
 sg13g2_dfrbp_1 _373_ (.CLK(net17),
    .RESET_B(net27),
    .D(net3),
    .Q_N(_157_),
    .Q(\u_top_module.u_i2s_rx_64x.lrclk_prev ));
 sg13g2_dfrbp_1 _374_ (.CLK(net17),
    .RESET_B(net27),
    .D(_040_),
    .Q_N(_156_),
    .Q(\u_top_module.i2s_data_L[8] ));
 sg13g2_dfrbp_1 _375_ (.CLK(net16),
    .RESET_B(net26),
    .D(_041_),
    .Q_N(_155_),
    .Q(\u_top_module.i2s_data_L[9] ));
 sg13g2_dfrbp_1 _376_ (.CLK(net16),
    .RESET_B(net26),
    .D(_042_),
    .Q_N(_154_),
    .Q(\u_top_module.i2s_data_L[10] ));
 sg13g2_dfrbp_1 _377_ (.CLK(net16),
    .RESET_B(net26),
    .D(_043_),
    .Q_N(_153_),
    .Q(\u_top_module.i2s_data_L[11] ));
 sg13g2_dfrbp_1 _378_ (.CLK(net13),
    .RESET_B(net23),
    .D(_044_),
    .Q_N(_152_),
    .Q(\u_top_module.i2s_data_L[12] ));
 sg13g2_dfrbp_1 _379_ (.CLK(net13),
    .RESET_B(net23),
    .D(_045_),
    .Q_N(_151_),
    .Q(\u_top_module.i2s_data_L[13] ));
 sg13g2_dfrbp_1 _380_ (.CLK(net11),
    .RESET_B(net21),
    .D(_046_),
    .Q_N(_150_),
    .Q(\u_top_module.i2s_data_L[14] ));
 sg13g2_dfrbp_1 _381_ (.CLK(net11),
    .RESET_B(net21),
    .D(_047_),
    .Q_N(_192_),
    .Q(\u_top_module.i2s_data_L[15] ));
 sg13g2_dfrbp_1 _382_ (.CLK(net18),
    .RESET_B(net28),
    .D(_000_),
    .Q_N(_193_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[0] ));
 sg13g2_dfrbp_1 _383_ (.CLK(net18),
    .RESET_B(net28),
    .D(_001_),
    .Q_N(_194_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[1] ));
 sg13g2_dfrbp_1 _384_ (.CLK(net18),
    .RESET_B(net28),
    .D(_002_),
    .Q_N(_195_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[2] ));
 sg13g2_dfrbp_1 _385_ (.CLK(net18),
    .RESET_B(net28),
    .D(_003_),
    .Q_N(_196_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[3] ));
 sg13g2_dfrbp_1 _386_ (.CLK(net18),
    .RESET_B(net28),
    .D(_004_),
    .Q_N(_197_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[4] ));
 sg13g2_dfrbp_1 _387_ (.CLK(net18),
    .RESET_B(net28),
    .D(_005_),
    .Q_N(_149_),
    .Q(\u_top_module.u_i2s_rx_64x.bit_count[5] ));
 sg13g2_dfrbp_1 _388_ (.CLK(net15),
    .RESET_B(net25),
    .D(_048_),
    .Q_N(_148_),
    .Q(\u_top_module.i2s_data_R[8] ));
 sg13g2_dfrbp_1 _389_ (.CLK(net15),
    .RESET_B(net25),
    .D(_049_),
    .Q_N(_147_),
    .Q(\u_top_module.i2s_data_R[9] ));
 sg13g2_dfrbp_1 _390_ (.CLK(net12),
    .RESET_B(net22),
    .D(_050_),
    .Q_N(_146_),
    .Q(\u_top_module.i2s_data_R[10] ));
 sg13g2_dfrbp_1 _391_ (.CLK(net12),
    .RESET_B(net22),
    .D(_051_),
    .Q_N(_145_),
    .Q(\u_top_module.i2s_data_R[11] ));
 sg13g2_dfrbp_1 _392_ (.CLK(net10),
    .RESET_B(net20),
    .D(_052_),
    .Q_N(_144_),
    .Q(\u_top_module.i2s_data_R[12] ));
 sg13g2_dfrbp_1 _393_ (.CLK(net10),
    .RESET_B(net20),
    .D(_053_),
    .Q_N(_143_),
    .Q(\u_top_module.i2s_data_R[13] ));
 sg13g2_dfrbp_1 _394_ (.CLK(net10),
    .RESET_B(net20),
    .D(_054_),
    .Q_N(_142_),
    .Q(\u_top_module.i2s_data_R[14] ));
 sg13g2_dfrbp_1 _395_ (.CLK(net10),
    .RESET_B(net20),
    .D(_055_),
    .Q_N(_141_),
    .Q(\u_top_module.i2s_data_R[15] ));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_31 (.L_LO(net31));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_32 (.L_LO(net32));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_33 (.L_LO(net33));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_34 (.L_LO(net34));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_35 (.L_LO(net35));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_36 (.L_LO(net36));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_37 (.L_LO(net37));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_38 (.L_LO(net38));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_39 (.L_LO(net39));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_40 (.L_LO(net40));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_41 (.L_LO(net41));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_42 (.L_LO(net42));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_43 (.L_LO(net43));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_44 (.L_LO(net44));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_45 (.L_LO(net45));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_46 (.L_LO(net46));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_47 (.L_LO(net47));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_48 (.L_LO(net48));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_49 (.L_LO(net49));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_50 (.L_LO(net50));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_51 (.L_LO(net51));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _418_ (.A(\u_top_module.left_channel ),
    .X(uo_out[0]));
 sg13g2_buf_1 _419_ (.A(\u_top_module.right_channel ),
    .X(uo_out[1]));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_4 fanout5 (.X(net5),
    .A(net6));
 sg13g2_buf_2 fanout6 (.A(net7),
    .X(net6));
 sg13g2_buf_4 fanout7 (.X(net7),
    .A(_138_));
 sg13g2_buf_4 fanout8 (.X(net8),
    .A(_100_));
 sg13g2_buf_4 fanout9 (.X(net9),
    .A(_099_));
 sg13g2_buf_2 fanout10 (.A(net14),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(net14),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(net14),
    .X(net12));
 sg13g2_buf_1 fanout13 (.A(net14),
    .X(net13));
 sg13g2_buf_1 fanout14 (.A(net2),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(net19),
    .X(net15));
 sg13g2_buf_1 fanout16 (.A(net19),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(net18),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(net19),
    .X(net18));
 sg13g2_buf_1 fanout19 (.A(net2),
    .X(net19));
 sg13g2_buf_4 fanout20 (.X(net20),
    .A(net24));
 sg13g2_buf_4 fanout21 (.X(net21),
    .A(net24));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(net24));
 sg13g2_buf_2 fanout23 (.A(net24),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(net1),
    .X(net24));
 sg13g2_buf_4 fanout25 (.X(net25),
    .A(net29));
 sg13g2_buf_2 fanout26 (.A(net29),
    .X(net26));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(net28));
 sg13g2_buf_4 fanout28 (.X(net28),
    .A(net29));
 sg13g2_buf_2 fanout29 (.A(net1),
    .X(net29));
 sg13g2_tielo tt_um_i2s_to_pwm_arghunter_30 (.L_LO(net30));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_241 ();
 sg13g2_decap_8 FILLER_24_248 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_8 FILLER_24_269 ();
 sg13g2_fill_1 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_297 ();
 sg13g2_decap_8 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_311 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_decap_8 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_8 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_fill_2 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_decap_4 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_4 FILLER_26_357 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_4 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_4 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_4 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_decap_4 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_294 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_339 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_227 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_4 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_4 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_215 ();
 sg13g2_decap_4 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_decap_8 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_decap_4 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_357 ();
 assign uio_oe[0] = net30;
 assign uio_oe[1] = net31;
 assign uio_oe[2] = net32;
 assign uio_oe[3] = net33;
 assign uio_oe[4] = net34;
 assign uio_oe[5] = net35;
 assign uio_oe[6] = net36;
 assign uio_oe[7] = net37;
 assign uio_out[0] = net38;
 assign uio_out[1] = net39;
 assign uio_out[2] = net40;
 assign uio_out[3] = net41;
 assign uio_out[4] = net42;
 assign uio_out[5] = net43;
 assign uio_out[6] = net44;
 assign uio_out[7] = net45;
 assign uo_out[2] = net46;
 assign uo_out[3] = net47;
 assign uo_out[4] = net48;
 assign uo_out[5] = net49;
 assign uo_out[6] = net50;
 assign uo_out[7] = net51;
endmodule
